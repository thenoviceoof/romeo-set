��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�ϗ7�#���H�����u�g[iˬ���t|�3���ҥ�ys�B�@Yq�"F}�\"QY����#�ڇ7�\ӷ��繟��1W�k���q�u ���{�m)RM�S|@�����ͣz��yʿG��O�Yg>�s$h_!��-~���=wx�=�M�����/�mb�K#�� ��1��W�i�{,?�EM�N�0�K
䧣�:39ok^�(��-���V�f���Sk�	����}ؖŸ�*����~������6l@ޱ����t����_.��±7�Eۨ[�ܐb\T�8�����"��!'���^C�he�K�Zw��J�;��E���a�BnB��lje8�i�U��^w�K�@ܚ��^<'�������������a}��a��W��S��!�P�:�ޓ��|=ǎO�k�σf&�_ K(yǦ�+F{v5�X�x!}e�y�D��"љn3]��6:�Ѳ=&:_��h�,�klf�es�4�=|��-�#3��r�E8m>�e7�{�~w���O3��{	 X�n���7��[��{d�mҫFG�6�ݝZ���4́���GF��yw�D��Օ��挹O����[�K6���L���ڹ�\Z'�
���lS}d}��w7�� ^$�j_��묡X<P�`��&X���xRq�y��G���R��B�}[�b50t��j�k\��Ju�a�V�ؒ���w�\%RF�Z�購�:*EO�GT+���,��B�/�9K�5J���t	���y"q��yǕR�<�]���>{�t�f�'z�(*��l�����'J|N�]�F����Yz�ȅy��/��)�B��
�vu`o9M5|�Z�e������gM"���C�W��f,�o�`��<��Xk�:�s#�T��/q�PC���k�!}5������j��b%׊a1-�b��\%猢��S������Ew�Z���UYwds�i��;�IT'q��z9}j��!/m�n��4�Z������ء�\��0d��>�fZ{�>�Q���}o�x�/=̪Y�I�s<T�y-���G���_�җ���2���5�g�$K�+�'y��wj�%��� ����s�ٸe�p{��V�$C����FQTX5��)w�"��c��Lg+Z�fvV@4�ZP�>l���
�U��������tAĪj�k��V����>lv�C�/8��M�jR0�:q����Tԅg%�L�:�����t}W�/vF�XȰu���*_=�Ҧ�/W �W�J��k2|�v����Q�o�2�l� �@��n�S&E����q;�Ǹ�(�b�?��&�pAM�� k;Eb���7��U�U�k�и}8�+9$��'����ݧa#{�~P�C@�u`�#����]�S�N{"C=l
�i��+*<�L�n�k��STA��s�%�X;�y��@����L����n��e���-�4���=���t�X�	���B�`�K�C���Ɍb��8!5te���i� �������9�E�y�w��ܺZz�
�5�_�w�.W%x���|�	
�Z�� /��x���f�-H>��|�)O�(�x��:E��&��Ͳ�Q����<>�E������B����
\�t΍��9��Ȟ��\���$�z`�� �1n@4/��e�P��$���u-��?�J�$?���Q�Mʕ��[��y��ن@0ha,��t�H���OD0�p�{O��M=f~-�G����(*��!m�Es'�#�A~�G���yk"�ї�����!A.���Qձ�&Yeis?ޖ`r4��9��7H�͚J9i�Ň�yʣ]��,�y��)�Wz1����?����Wt����� ���� �mT��"�\<��o�����D���^ϝe�x鞾�F̂���ˁ��ͪ΢:yz���Jc
��CN�!=�,�]$a�����Ù���2���rTc���Z�=HZ�$�Z��^T�{)�ȧ���_ׇ߹k ݧ �dظ�z����*����D��٥=ɬWb�	օ�����^���Ar�pLPH�7��G(�.O�]\��Snf�ǯy��(za:e�^������.�Ƭ�r}�GMP�s �Ǭ�����O�x����Y�T��3��`��3h�s:����\2�d�;n-�q8���FW��>3�|o�
|�ÿ��F4I����[Lb�8��9'�Yj�l���[T��i�V��p���eƤ��h�9���`=����[Pf��c���#����4�7����Y.@�ݧ��{��Q�MDm��D������C��2��]�4���vK��B����s�6'.s;�Z�U�e9J�:9�7��@T�_��ꐜ�M�x��>�`�� ���"�k�(V�я�����5��GS����ׂk�M���I	ǳS��Q�N��P�ĜF�GA���Wy�j-���D�k�*��M����ՒJ	�q���Y۩>q�S���R�(Em�F��\���-�h���Pj	M4oı����DN�����(,�,�|��SO!A�5��.��2�ɉz�	�K���q�'�=[ʭ|LX��Q�h;vn�S;̝�Є�%/o�f?*���[�B*�z��K4��)�D�gz��+.ݕ��c��%�V{X,,7+M�0cc��;L�W���zo��ϖQ���"�L7�k��1�鲾ě@�uo#]��` �00�v�3)��e�o�g9Д�(�e�$��5�z�m�7*'��
�.�J��ly�L:,ۨWu0B٤����?��RĘB+%yY�|�Q@������¯C>�<卓���<X�dI���I:�!�r�4+#(lpؒ&1���эb_�+V"������a!!�h4�B��PS@ {4�i.����eG�\�w9v��<��pp풥�OYY�0������Co�gFFp�[�|o�s��u��-W/�Hx�o3p�+F�;Lг6]6b��$�^W(�,ބ$���(�?�g&kyt_�e���s5���VE����{l8ݎ��Z�x�'8�^+��Wl8˧N�]v�Xѡ�t �m\K ���a����)\�$J{�[�=�4��h�}�iy2Z��TDy2@��k�N0��~���qt�x)�{��N<��LW`��uT�*���(�;�)��)���@N{��'zoT)G� B|e�eH\�(8���@�,�V�6����r��_8K�E:��&w �aeC�&f.f\*������2�e��C����<���
0�?��u\kYA^M��*��i^�X	��0]Zs��))�z	��l��8k�aNe2��i��3V5��]��zv��� f�\��$��Oƺ����Ni.�q-�Ӭ#��X�	O6�<�)��c�Xͱ�3��X�Qw���8RJ�x�(��xsC�-�
;Տ����px��'lHR
��Z��{|�{�1,
 �e7ų��	f��������~�GPV�S5U��0���(�ẗx4��������W��H;�*����j�;��������f�������D�Q�H�Nڡ��gT�Aw75��7�:�C�X��4�>�<%�i�Z;n5�VJU}!�0��zu3���ky��`0��M��
��j����eqw��T�xvB�c�1EzhMP]0X�X
"4p@HHW$�ik\9��D�{����i��Ԉ<�2M�v���,�@-q�%v2���,�=��埱�lѕ#��
%Z˓u��O�
�q�:0m����K�Pu�!0�;���j�\�Kyv�k[�0z�GN����ժ��R�Y8-&����i�]d���� ǹҷ��c�&�qO�&o.F�Eg�=A#%0`�Jn��U5�I!�d�l�J�J���V2Ylie�K��:_BĘ���;�����.B�|d��`�g�- {�y�Jl��L��&r�6 x�M"�p{�[�{Wc�=�!�ٓ.ۓۋ_��I[n^�� L^�
��2���I�R@쒬���H�n}��ఉ�y�fÅ	���>�,r�-�-^�<1�L��$��h˰���L��X�ibI/�K�J��jXc�n��w<�A�J��ȅ?����N�ݤ�z��5H���ߺ�=x��S�ˉVH�x���Ր����p��O(#	�ӽݸ�� '���⩊<0�v�o����V*��Kr-�I
�w		Ŗ��i��|����9|��N�3�
(=��0Sh�@˔��f��Un�6�V5Վx����o��B<�99?P.��/ H����gY#0�<	��� ��+PZ�E�V��)�J
��s���.�N�ΙyŽV���_I��O,��`�'��<|��YЗ�[�QҨZe�T��B�0\�R�:�&�>�B�Nݠ�,ʝ����/��� u�=A����#��d�
z�U�x�5����T��4�sK���m��E5�rfcg9bx���ʶN��V!�Y������)#-D�+)��9D�$���+iV�9�SaP�	�p�~>r�o���n17�7RRZA77e�)*D���˄ߣ�d�f��������)�%��< J�v��)4nO�D�Q�)�wDX5�@a��=�;�7��a_w�OR�zw�r睟�;1�?���17�0F4OaQ���܎��Fk��bp�k��o{��u�������?z��dl�+�H[m��5��xg�#3&4}����J4�
(U��Q�-���3x�T&4H��(����|"��Z.��
���hN���Llk~n�q�A��1��x��Gޓ����bt$���pԸ�P��K4Ķp����w�Kf,8{k�dA�i�p7��֩�i�~}�G�d�Jn/��1?>�n,�i~�n�sh��D���g)O5X��u$+�f���V�z���\(xL՝\�GaIrE/`;�&���m.�7
�\��y4�Ie^S��/u���V1���?���B�e[ '��{��SB� *6���k��� KR����z�����h��g�x�ǭ�ʧ�Č����J;)s'W=w���z�9Ich)=�_�#8�{���\����=�/�`/����ԂapQ�����X�+�^j���`0H�t^͋�Z���u�R�Nl)$�^�w�*<�xG����.����Y���Qp�wu�y`����R�Zj��@�ery���y��	ܠ���w���$�]u`1�f���pd]ӏj��u��&�fU��¤��7��K�>^FA@gp�
��J��N�l��[P��k�Q�����Fy���Un#g	��g��'�mO*��P���N���1�>W��c��l����Nֈ�=��k���6�fsm;�\o��m$hjAW~$��a��o��`�@�c�=7»9u�{^��%�ؤv�F|{c�;ǉ+ac B�f�R�3�g�S��J�Z8�)р���F�OA'y�[��⫖%
�L �0�}żА�f���,^���kи�>l���Hf����j��G%�=�ܣr����dYD}q �y��Hf�
x����F���8#�B�R����s�[�m�Ow�C��"���F)�ޜ6iP��k��ӹ�z����T�;�o�Q���×HE���n� ���z�f��?:N�s��(�j��W*s��u�f8}�U�K5�#a�5+��V�bKI�R�K�rQ�a|�U]��xq�����n���]&%�\�/�a^�:�3Jkc�'l�n��ǎ�5(0Hש-�u��J�z{���@�1Wӆ�̀��������VCQ	K%kl�b.�<�Sx����c�Ü�B�w�1ڙb;u��Ʊ�������50X�hr2�G:�����JI�'�IO�V;Q)+�V���.��wh��.4*�gH:	�(7-��[X�DT�L���j,ӏ[���e8�'xd�O���*���Yrnx(������x&,K�<���d�SU�ߗ��J	�7��J?H�ڒ�@�f�p�"ћT�#%�E/}�K����>:E�����k�R.��Q/��7���%�ʪ�b��|�/1�b���谕�TS���~���*�5GKf�/qk����F��TkF'��ReY�KmVv/����-B2 �`��j$����M�FGC�`Y����EB�I�e����P]N/:��9�_�����N.��s��s���4]�aI�5�
�l��N�M��5����W�!�]f[���h1Ħ	��Ń�_ZX�l�է賁�U^Y�E2|��lƉ��^[)�G�����8�%2�0X�D�t��¿?B�O�7���ū̠�8�N�"8�;-�j!����Wk�}/����ȳr�6�(�e�}T��2�U�P+@ސ�ӆ���AϮ�R7D�D�/+��oC�1�U�#�i��_p�4�3��G%�]#��NwN�zY��Vۧth���������TL�`�3g�;�e�a�@L?���t�mOWX�p�s:�V����a�����C�!_�I�w�)���a�������xُ�+����R ��(T�ierUc�4���t+!��cO0=n��+�CDp�!}g0��I���jH �A;:.4bYv��#�w�O���c9�@	�K�5���Z��
�$.��c�+���cr�3d��$Ч��ˬ$�G�-��n�%L������Fdi2������t�H�y�,���v �$�=Ͻ���9��[��r��5��9�J>��T,��X����ʟ��EQ��)|,��C�]8�����y|dާ*��D~����#Un+~.�$�x#b��v4����v�=�Ohيr_���1敾W�	������p��1�t�.4æ�e4~��"8/V������|*������贼�((@��]{Z��H�� ���\�s�w�G���q't����[!`t,wNV�8㾽�-_q3��hD�6H���%fv-��4���a8��5�N:�)�[���_l��F�yXX�������+��x&`,��Z�`��7?g�/b�ɀ �9����/���o.1Ʒv4k=��z����Xn���0�Y�4!���A�!���mK�{��FE��Ww8��qeVd(�%J¹���0��ܹ��;L#0ݱ=���]P�j��"]��i�CC�&�GZ�VY�+#C�a�@E@���2�� -"'�xf��s��6�mY2.	��P/�G��$s|��AU.�M=��+p«3TF�Y�@t,�Qb
��5�Xj|�*8��n4�]��ii�l��Y6,c��1\���&�����k���e1�m�<������T�=:�#��Uy:2�� a�C6�0�gܛ�q,Ix����Z����-�e�JB� jnJ`��~�1�q��ڀ���2�j�Q:�@?b��1��;��,x&b '�8?�`S#��B����&��iB�]@�L�#�/o[�oI�
�:�4��o�ͬ)�K���@��
Nf<$���m/!�"�׏��3� �����T��Ƒ��=��y�-�r�1! ��1ix_����v�3BR7���I�]��)PS�ҧ��f_kA����Q?m�������hc���P�z%��,~k���w�Ͷ��Ξa�Q��ܪr/�t�EuP���6�f�������a�����W_�J@KL�9�`�#��-疩/bl�FW!1�����*�����wZ�)��f���ԃ��J�A�.�h�@C'�����*�T�~��"=��rL' �vC���I�{�- ���&!K(�.�s�����P-��4�Fo���E��w�s� ⢽]���-\O'�߹d�U�	�jH��ԝf4�;rG*D�_6������~P!Z?�;wА�T�T8]�_�>�)M�����tXz=�{���4��rץ(i]�v��Lhϟ�fś!Y�K��m#�/���~�J�	����*�o#\�H�!>3}-����Nl��M�m�__o�`���R�5���R�e���'5Q�Yo����Ø��ԡH��U��t2�o�	�		�*��c�lxe �WEmK��z2��347Ԛi���䩰��bl�Y~��f��Wؾs�ڝ�&Ϳ�	���~'k�gC'���&7K� ���œ9!�;�Ш�"�9����SrEƷ�������Wo0�f%l"�A�M������Nx�9�~#�-Oy�e������Yʛ�=P�[\�o���)ga.�� C��߶gk	w\���w9~l��z5Y�ڻ(�`��,�U����<����kd<"�Fk����i 2�*߻�����m�i����*`��Zɕ��:+�5R/�,M�lb�O��.�� �s��ۓ�e���sY�j�w�P�ku�bm�D|�G'���I�;{���n��&�&��{��4fk+�[���0#��u��%�YǷ���D���ޜꤲ\yjK��~Ɯ��1l���
������i49��\odf��'����$�ۤH;�R���}	]G���T��uZZ�{@ߒOzQ�TY����!�z����ī�jL�n��m����4�sEu�Q�-�	�,5ёZ��C�*uɇ��?'�G�;Ek���ʣ�[��f�;l*�д�#�斡�{��߂��=���"�z��KR��r8]��D7X(�ﴥ��"K��$��|Ao&��v�����75jV,Nh\dΞ�� �I�%h-��C���Yy�1q*j���qN��~������]gG�L�m"k>�����:\���٦' �O\����E���׊���;��;^&ժ�k�P@�·3�z�eȲ-�N \�|�}"�h�e0�����'M�`�x�R�U�"��6�ܳ��ou�ȋ%C��������I�<R��������N�@��J�ٶ�٬�u>;����x��ýCۦ�25�N�S6� �dS�b�y������c���U>Y[|����W�D�;c)f���YY��ELtN]�wg]���.T�c }�f��$tեn�����Y?W�NO��8�w+~]_�*���2�x�e�bq���F��	��bp�$��=5-譖I-3��Bj�?"!�v���A�Q��	��%��c{>o��!�Vޤ����j����b`�P�w}� �dJs)׍Ci�Ej��$��wk���\�
����.8ɲTݑ�^�h��L��?�F��a.dZZ�d�f'gF�7d^ h�ۈ0�I�汓�=�|��^kla+�O���N
�+�S�>zxM��d��U�P��{C�L�Bv�v4̿����q���\��k�G\)/ Q砷D�ǌ}��I���1�&�����ZtN�*�H>d	�3l�V�@��`]����Q��YU��1�#K��?N&�=5��|��ž�%1&���u�)�T�ڞ��p}8��o�����y#�)�����5�5:�'�ũQי&�'��5h��{ֈ��|Q��8
�i �'Om��CK�w��=Vlos�n���a4H&+ؕ�n�{g�|VW�W���LÌ\�Ne%΄�X��h/b-�k	�joz�.�Sn�k��!Ƭ��6���Z����5�;��x@�~Q�˙�ɿ%��='�3�{#���{jᚱ���r�f`��_��+5�&Q����� +M�/���g�@�񡰧�Q�̽U��ꜿC���;��T]�a%S����y�e�e����5:	����b�m�.��Z�5�;;�a��EZE�o�N� iީt�������V^7d�pr���Rʉ5�R����W�5C	�R�y�y<(�wH�o?����.�Qp�DK�}&HG��38\h��/o�\��w<h���Dd;_�cїlX��D�^$/�ۭ̐ߠ��E��?��j�Yz��OE¡՟!U��@S}�G4zj�m=tr��0����ۼ H
�hՄ�OZM��B+���S�(��<��E��>�J�5D�k�0otN�T��Q��Gh�6���^ѷ����3��p#j/�O���� 7���n؈QXܢ���w�u��c�AX�^O~��'^�I3h]�����4sώL!Vr�7��	�g<8a���$i;�
�{0�p*�}�vv��#q�9y}֎6b���l'�Ә�D�Y�EfX�@������5p�����s~�������c�?�4��Y����?��*�s�PK2 �x���x���w��)���X��\��f��K��""�Cx���y�$~�BRvݧY������*�xUhnrY*��Z�U!�%X{�
��T�F�H^툉��s�
ncX�춼�7��\��w�v��$�T�)��w����yp����ICXuu��H�f�:�ִ���<�*Ӭ����9���
���B�ž _�ݥ����HH(C^�#-;��KZ�%�ǐ�D>���?���-9�9<Ԥ��u����_��E�[ꇘa5/Ia�f ����"z^��}H�`첒-�k�)�u:٬9�8U�6�ݎ�~A�E���D��z�h���S��b�W���A��n����*A�%�sf^ �2+�{�by��uַ�#xt�~���*� eT����N�d�����ms��+c���
[�*q�s�*��d,�b�M����͕��7�h���e���{=#�����]��0�I�q8n��h<�P����Q�O���,@4/lS�PZ�ar�&����ƕ�X�=��-P<����&�c^��d��;�`��Ve�^�5����'"'؅�X)(S&�z���J��<�vT��`�'�q�Q�a��%��6Ϳx0��hȡ�pO *u�-��Q��	?C����u����E�C���O{R>�;�Vo��]�J�~��5�:f~. ��r��ͥ|s��9T#A�g����.�����~r������96�7SROT��R��g ��KԞw���G7ߣ�6�u�tn:&��6��|l����K"�(�&�|� K�'���{|f���-ؚWy!��8��?۹�K�\�U���b	��v
�l�������WWh���x�H�����es��b���#!{%����*�-}�{NwK��RۿiX/�Z͜p1�o��nma��-0���;+��t�a�j��4Մ��i4�i��X�rp"���W����S��d椗���%�?�g/�9�c�p��x�4�w
�7@Gpr�P������o��epvRK���J��Ҥ?r����''x+s	|m��;�v���> ���IYH겆���6k���L�O���3 �^a�%y��P��+;��u��yg�`��+k\�������p�=*y�j��r�
��C#�<�^r����V�dv�r��X����!����сj-�[���.�./��T���;^����/A���0�r����3����q#��e+��V��E�L��~� ��h���}��H�]{&k>*��l0�Ne#�b�)�ҕ�8	A]�{썌��*�ʠ<�.K�fVe�fS��*63�5Ӟy�4��?�R�9ǟj�1��_���Cb ���PF4��@T8�e�����1߲H��W��gY{���)�����і+ח�lgk2�������6wq���)��v.����Y��Q� �>	�&q�`�����S������g�e��&����&6^ོ���ir�.(����r6uJbF��\oGo�
�bE1P��/�;M��6-a|�A��T�('Q!
�T�v-�S!�̈́_�9��b9->oM|c"�Y\Tn����df��+�*����-�:ni��jM�7座_��B�^�u"ͩ ��%4�s�I�s�z������z��c[�4��˦��7����+�`���S���#g�~�`�@:�s1�g2�p���[���k�$�V�ɲ+x<h&�#��fp2�A�A�7]����Y�W/%G�I�1W
��\�s.�Tu�t~kdW��~�-����Mh����=ܟl��QV�51�SX�,�]�fHWU9�h���oa�՚ ���
J��t�!�;H��~}i7�<�t�0c%D�>��q&;x�F�d�f�n�
�w�Iȯ��i7D�R� 3�p&�%��F�m>�E+n��FI�eϒ��GT�8F]?�e���rV�"�6I�W'ĉ�&dMP�B�5���5��:~��A�=j�2F�(Ø-�կ�?�|e�#2��W�nE���I���C���Q,�oe�շ�)b�!B^�h�km���L���(>���Nk��ۉ�b�Z�/e�TE2�Ͳe��6`dv8��k�����Q��j��Ks�E��q�W�Uc�"�XYz�w%%#쬏6Tx�����
���L�� $��>�;�ѻ�������ϧoe*���S�"�ǩ�E��y�8$
P7!,�E�����
�!+�Q9�c�*�@o�D�L�߫Q�Es�M���<�n��7�F�t��A0kI�Pg5����0!ͦp~i1�lՉ��C� !w< �� �}�����o���v�ҏC(;������`4wϪ^��An��m0�� �=?:1���e�-�9�mՄ�CL��g�e9�>Bv/82,�xgS	���@ ��Ly�,�����;�L'bzϦn!�g�wG^�f,c�N�/��	��N<@�k�.s�\���B�~�7�)c�GM6J�qW�]j޽�Y��Vn�ږη=yL����o�]�S6ĺX��c/a���(��.�t]т�_P�G�<c]��/�L� ?�����"���N�upwMٔ+	��fD��N��e�L˥m.��`�9Z�۰C42�_
J��B/��v�XU��L����^r�uv�r֪�-Z��v4����)r�ۣ�:4�����?\��eD�6"�4�̠-�����!V�Ug��y�9r�ujpXϽ��a�sP.h�JS��T�]��B��v�r�.ѕ?��m�'O��j�S9̌v���4������6�X�8׌��H�"p6yYF�q<�����Oׄ+��nZo��h�!�[.��b�E����`E��K6��n(N�n튱���2�P���c�'��������V n�
�]>�e��˓����O���fP�nN�Vgc���w���h�QBm�W�N��T�Z�wCX�����W�#I��W�Z�i���^�,.W��(A�C�*A�,#�>aϵa!�L>ۅG;f�=+*(����]����ϫRV�Ƭ�Ǟq{�gY�������<! d���+3�>��[�)m?��N��z�QLZ[[(M��w�ʱ�\�6�b"�޹|1Ȼ���FV���T�DID�p$+aoc�P:�t͉n�����a� 2�G�ż�����O9�=��I���T�1�S�Žp���rZ�0Q��NK7�2���N��vD�ێ�z��$2z�T�F�b��@�@o�;�I]��y���=�3�_������yd~;"�<����Y��P z�b��8Y��l7>���ϧ{�(+�q�Y/~Xt����$�.��{Ǌ۲F��m�4%Ѯ�����*	@U�"���?j֞Y�+V;|��VH���T���d*���S~k����_>��������#e�	wC_1�&�ў�!���~͹���[�k��2h��{h�UwW�>|:0�nȈ�FGe͒�%��'�����e|����b�]F7�Np,r����5Fd�!2|?�����`�i>VMT��X1)E�������p�c��*��\rfݽ�c�QsmY��J6	�q�׋V�fK%r���h��ћ���ޣI;�b@A�S+�Rqb����o_"C�������W�J�/����59t��Gd������b�<&�9�ߤ�$�N��5Z}�����U���W1�ӽ.~�3
?t"���H����T�s|��Y6�d�����N�q���bN����D��ŖL%��b���>�T�ٽ�4%<C�>W��f��`s#^���@I��dl-|�׼��0��&��K=*�G�C�kX��T2�k�RMI��Z|�����ݍ�j����6T3�����^f�p� ����~�U���:7;�f�S'ep��^�N�D�Bs�����k��%d�laB��O���*�����x㚶�wbj~�G7a���� ��)I�?,?3р�%U(M���%��6��!$e�"�:sUX;^2=�x�h��frș�����>	e�~]�U�1���\�:�2R���A;]�%�*o��:���N��Zy�T�����`�=?���Sq��JW�O		{�- w/#�S�H�P��/C����?R3|���й�zmO[똿dkfS�!�޳<g�V�a����t�N�V-� �eȪX%b�(�)#DoN}T�xNW��52Ӭ�܉�J�-���3��'���r]�DyGC&�����n��Hk�9O�[��#�����̣�%�w�C�+x�pi>S�ȑ����������~�'��+��Cv�m��IX�)n��R�"����Ƶ�S���)]G����[����IF��Ѿ
L̺�Ke�J��,�i�APV������K����a����D}h����S0EAKTCK�]��j��?�sd��A<C	åCW���NE��6	aΛ���./>��k񊯚p���&�?G�sO!,>W{��v��w=��ZJSz!*3��1*��Q���҃�0�ڐQ��m�Hΐ�3-�Mx��\�G�eQy~��#X�4ϟV��%YH�7a�0�7P�\`Q?��5V<E�*�xН��r�Z��[9nv��Z�Fb���e��8�hd�����+;:P��	�'�O����J/�e����ޮP��w�t>��k��	�����=��ɞ�*��H;`��Ǹ�*J���b�*0ko�7�W0^քىSKVzה+n�����F��tk�wh�e)Δ�m��ʝ
�Vv�k	�����
R�*3\<jm�P �pX�l��m�bڪ��J��^��������6wq��:"�TQ��(k��A�m�VlD�o�7g9�Ri.kD�����Q HdP�/p�Gw�PXTEB�&��/�dGCn�������u
�63��T��� �����{�f !;t���g������R�8�6�a��k����]��ܭѴN2�gt�6A?��YK-�$���@^}<��m9(��#�����cy!$o5:DC�ev�B����F0�'�s�1HG�	1o���Г�X����r��>��.�IPY���5�� ΃�8�\�A
��0:������_mbE�nM?C�J
����Dm��e7sAs��s�sfR]�!���F/�C�8�ܻ��)ҝ�?�s[C��x��TvBN�+.�J�ǋ��n��nkK;L,,�{L�i�i\}pB�T�B�S�}���-�M�*����0��#:�j˕! @��Me@�	9w3��`�a��ޯ���B#ߴoҵ�b~������Z� F,�ŅҾ��Ē����q��kJ���_�)��Vv�ת?
_t=�2t�1OoH��'(+l��^��`+��7��RΈ�0��7&U�o_?��'?�v�0���\O�!�<raa����n��"�_8�c�Ժ�u%~;��Q���kD��K�%V��E��^��_�W-��:lUđ���3,T{�V�Ou^/YK�x�gD��d��"3�HMkX�?�|��äje�=��;9��;��h#�f4���k�u(e���h����g�ȍ~�����e����᳸�hS�0�L�Ӵ
�R_��PE�b4�C{�99�ky*ɮ3��*���±�K���7�G�dv6��>��ہ�l�'�_cҌ�� 60��ZR�@n�j�m���꼙9+�5�*��E�h�'.�CC�6��f�|1�Ǒسp�oȬOL�N����.%�Fn�j�=cs����[���S܇��S��
��v����|��o:4i�
�X�<g],�{)�G�!��g�uV�3�ѩk���ٍ���D��]j���ғ
xL��;#�i}NxR߳��*5:I�Ȫ���� n1��gy�7��FW�tԩ�AՁ�wh�ěҬ� �"\k��#o��]���"��UP�3a]�,�ү�}@�I��RJ<�#�1����� ����դ�@o1#߻����ܠ�h}�o���3>�r�ks<�G�r��<�@�	#���
�����D�J�򘩴h�6��'��ȏ�sе��_Ri��%c�(��K�O"*AR3ϕ���)1�L z��l��~�Fu?���@Y I��<ʄ�a�'�͐����1@�|;���gw}�����X�7��)��1�9|�u\���-�4�^���	�A��]��m���l\�Nc�A�Ãg���uk��8⿈=��>�� �ܟ!EM���j����K�,��ߕ��"�,4��3�o, 3k���b諽sN�E~$6���>�b{��lɞ�����`��Z,���gB%�&lX���� ���E.��覸�ߘ_�e?&�]�� E�pS�˿Q#䔬���WUX!]�v���LIw&�,�7�u����ͯzU��6��Ȓ�[�'REd�\5Д�dϨH�H��, d7Rf�>�c�7�<o�\$<0ܪ���_9�h�q�IA�Y��*��o�l��eB�M�?̅���c4�D��PE��x�tDA����W��H�[D�ޥ���Q�>����\n8�z�!}���@�#n(�N�N�������\�ך���<���%���3��?m]�QM1bW�����d���xL��vnYs���;�n�:����,�P��TZ�e!��#�;t
��꤭��vf;� �=e+�&N��ߺ��QY�D:��-�p8v|I��N��˭�7i^ݱ>Vf���j���,�E�u��� {�N���pOVb:�2���czhl|��YpE��+�DG�����3��[#����*5�f�'�fl�d��YZ<ȧ�z�͸��q�3k���mg��!��!NC��/��9�����F�>w��Yғ9�={�l��,���Q��Ϛ���wޓҭgDP�����1�����V�1M-0��^�e��/�:�HZ��beQ#�(���ǧ�Π�i���f��垣��	�P{�B���9�('�"O@9qX��7�� �W�,�M� ����g5�I��r��Y������٤x�P�[��
&�h���ә�bU���;���HoHg�į(�W�c�#����`1�{�� �r�̺D#9{��<������"����Z&���r�>	����M<a��}}7xh.C����b[;k���3釮�mԓ��aL҅����ԯ%\������n�9v�F$9�56�n�dY�sq_SCOw�UY��?� ��T>��\����F�����tE�|������a��N}�}i��&3�Oz��AY7A�Ӕ�/���f~�&����2��N-�H;�(��IÙ�!t��Uؓ�{M���hM����e����ʙJ<�m����3;�H��
R�+̇
��??�̵?�ߒ�/��n�:]�9��h�� �O�p�l�V���E��^�]�mʨc#��+1j6p���S�"|G8#jf#�ԄD�R�F��x��d�;�ɭ����v5+�z����Nk���fZ-۶��H�6�O�J����V��[Ja�q��3��e��_�����"� �[�:��|��?D�D�[���=��|��:�0G],�B�t���n��M��v~̮��G`WnHY�i��О'\g?�! )ίR�k |㑶ё�9��<E����?��Or� 0�T~y ���i�Y�R/dy<Z����j�{U`(�W)ǴGv�RW~�ǅ"�Ѣ�*����R�e��n���M���^�Fo\7X����y���KN��Д�Z�
L.�7�a���ڟ4 O��G\
��{��7,�u��	z^S���O��I/�w)[���5�sZR���c�̚�C9ק�ք���ҡI4!��!��D��7�Ɂ����-�2�]䶙��Ə>�~)f���KU����8�[-�ЃY��� ��������$����f�W�8�p���m<_�G�[7�A��P{O.|�~��#��ik�����bʨ��Z��T���N-ՃJ��U���@�CV�-�mP����yU���$���,A�Cl���yd&�'L��=^�Z���ħ�G&.h�	4�ۍ݌{��z��0�f����*գ#	�>��c�sP��
O�s�F�����R�s�����ܡK���b��!��r1�D@�L^ɔ�7k?�#�N-��|܉��]���(ғ42�y�T".�;�"E:���3���܂yŃ�ό�Rۆ��s^�}���3T��
�uG�����_~�p0�n*�ɔ��pl�K�R���`�H �gT�����	@���*E ܇���2��{"s:��~�}V��?6�u�AKW�{@���Xv�7
AivEQ"��B��T������I�I��]'+a	�L#����U3c��Nd�|?Aw*�E_�o��F�A(]7�GY�#��]���U�:�v��.K�d�1�@G�ԥ�9~���H�G����]f�T��r�O�3���O�����%{BU��ղq.�&K	��v3c��\Rw�fH��b�e��Z0v,�l��G cP�K��N���<��:z��
�Fj�!�r�(
��;p�S��D���x����k/��fn��8���5��\��Mv�_e��sF��\SM�r�X���1j�k������*���=�N�,B>�:�5�欏��1��Ep��۠y) [��(�:�O�t X��_z�%;~+
����%�F����y��A__k�cqm#v�c�	C��!�8��}x��ܧ�����%��V����cʲ�y�/�����nGƀ@m&+��ے��7j`���QH~$"�_��UD2m��e(I����"����he/�JC�5ߙ|+��S��L%,Ĳ�	��v���H>H���|I6��|Q�Y�)DTd��ĭ}Y,#~���2�櫣�VXp���U��!%Q�L�\�pa�U�p�#*Ue���sx7���$�C�r8?M��)��X�<�J)]����������\��8ȻBվk� LM�%ߣk��h��Q�i='Q	�b���s����*Wo�R]í�j��܍q�(:�Q�	(���c}��1�*�|�&�A@����T4�i���l�����j>�o��L��|��b�����r��v���� �~}�>��yL��C��SiO"QOӛ����ţ��E`�:��_2�|���k"�+g>W4(-�A��1�%�pM�uן�X
��dC#�ϖ�&�S��0������{���5
���FSE\6pg��Y~ Vxï����Ȭ ��H!��{R�5���]G_����%%7ɯ
���S$�s����/�/ȟXw����P�x����6^R��p�#�g�<��p�fc�]�f3����4x8nW{+ X1�"	��Y-��2]��Pĩ��n�)*�f��@}��;Y"L:��kj0F(�%���Q*��}�Ñt>+L��dw��hB�.�xEH�h��e�D'�CRU$�p:�^I� ʑS�7������%C�@e�LطS3�f�Q-�ρ!��!��#C �o&�R�=������r��5k��^��?H�ȝ)�$0���o� �(���J1���N&��� �`.���H,�~����q
�K�S=��FW6F+�C`T�$t���	!`�0��@�\���$�,���:;D,&;�@,��!h���ޕb0<lO�7�s�����T����zx��{��C��z�I����%䤇1Ek�1��aw�SWm�|�S���Iv?�����
)����7Kα���و���=�
��k�#T����e(iR|_9��P�Ng�.��+:��g/-����u�;�'C���=�[����k�Ơ��S�S�'����[��K�CxB�G�TX�K���³̭�`:�V,���^��*d-Y�yD�s7����l@ �#�m4V���9�{铌�]����j�o����u7�I/��4�q�*5��b���r�k�i��L�����ܔ�WV�l�J��Ƚg�\\�'Hn��Ѫ8-�]�����5^��o������.x�*���0�zof��6�XoQ��U��f������6� [8J���9"v���lCe����A�97Ɲ�и�u���I<=��	�G��O��f��'���)�ٯb�R�SO3;���ެs��KE���oW���v��p�.�J\W��m���h�N�� 9X�71g�d@"��<\+�=(�2�}���~�|#ub+!�i��_t�������K�2�>.pu�C�L�*�w���"b�>�M=�0:��3��3��4HdU�!?x������X�G�oR�zҳ0���5Ĥ�P���#R�q��
9��������#i���l#]�� �NM���
ڦ?#j�>�	��'�= (��*�6����;�D��!�����:U�Q�ZGm���c؜JTm&h`��м1����y�69���&ȜV�a�ʨ�`@�V��{	}wD���6��.1�;W^Z���l���-�����"w p��d��4�3��P�߅e�x'���q��[�
<WAy�5x}�]oVf� �_$W�=^G�"�6C���������<O�| �\�8%������0�|�9 ����	�I��E���+�9(�
� `���i�XB�B��cb�[���HX����<�]�� J�zYr��6^��UX�ށ9�G��j�Ke)���eŊ0VA���&X�
R�I��,X�Ϭ&���iK��o���S��� $!�o�'�͠X~�͎m�����&=��P�2�ۙ̓�ݔ�t������ﭦ���{���a:����N�]�m�Գw��~�������{��i��6}����񛕎��	 ��1Rf��Sgyb*?"��]�k#6�Ɩ���m8��O�b��T�����Y�L��)���~�vu���Y�7��CByO����9420�Ϙ[��ߩ����ռG=���Ϲ��Ph��3Uz�'���̪���`(N����'��:����DJٝ�k0��ju�����RP
u�����Ԛ��|��7=zCJ�c���eOb=	�.����U��������ϡ|�7,�Ss��Ss���#�7���������kL�;B[���2՝�0V�m�\8x��\���J�E�l��i����$0HLCt,��#[�YvE�.�!f�J���]��H���m��D���ٌ�v��&���d6�P��>����Z3%(�2��ܢ���}@�q1@I	�QnW���A���6�4+����d���T[[ycJ2�z�-�W�V�� NU�jL�&Է���l���j+i�#��)Sa��_��m�N���]���7��=6-P0-�@<��a�z��3�݋�D�]t�S^?ye:�/�V�������Vt�d�ݥ�E{�����"�-�ηsqw��t�W����'��D���7�Ή��@u��*߅t�Q}],��qB����#��߭*7��J^YR\ů���,7���@(E��8k&\m�+�؃�^�f�5�2��G
���i�v���}�}f��hR#��i�	�Q��n(��l��կY�*�e��Rn״�u]*P�l�����%*�C�8��쓤���?����s;�;��.!��t���N
�ֵ�2�teSX�Y�pcP��y=��zF����O4*R+��;�z��?�|����o<bM��}vnh��J灶SO�������hM��`�!����4e��:�&gq�F�b��P^�Gb�h�|5�ې�dY��S��4C߹%��/��OU��8���������OA�%�5��7���� .<R]�Gi��Z�$؛'�w��^�����eh�jm��r���n� ���")h���t��9��S:=�Ͳ��x|N]p���rb҉��\�AN�nc�0������/t�G�8�G�����i�p�	~?	u�^���}�<X��3��ݲ��o�8g#E��X(цdG}���/��1�>gAPE�j{���},'�R���订C�؋�X���a�;-�_o���n���1H���/(��2�LU�\�q���Ps4�XT�o0G>�sl��^����v�^�թ,,�V+ȓ�Ӯ�k�D�K����!���^�ťjj��j��h�c�ŝ�����]��:�(�sy��n!K��LPn>����8m,$��2��T�Z�8'�0�t�Я	���Ѐ_a�v	�?R���H���V1�_��lV;�YO���%��J�=n��0�o ����s'2�/����~�}dL��o
��cjak~��!T�1�\(������a|������0�8��q�?p�m�N$��Y��s/W�֤�n�9nJo�ȩ��;
+�lPxg�E)d�JfÛ7Xa�������ǭ�HFx��	,?�+܌���Ǻ���u���z��� �����+ݭp�Ț��E�6wg�
�ٻ9+,{ "a�$�PF	�f�]>�	�>���"W�+�]fr���At���)���Α�<&��34TS��o>�g�L�ݏv|��"S�!���Zv�/������`�
F��--�����e�����M���#�pl:ƶq=���_�Ǟ6�1'J��Oq21������w��If]3������rx�~�`��{S�����N]Kh��f:�pR�#֟���;�z:Q�2Ō��!��_$�v3� �X���I��/��j<�_(Ϟ<�o$U��tg~�<��]@^Y��<_�]��e�xz~%C0�p!���p�1�FnD��@ߠ�p��YTb^�AS��d���"m� ���r�6m\Q�S��q�s�n�'��('�e����b?�¢)�H+�U�A{U�,�.i�k<i6O�R����G�b���1?X��R��[��YF�YX�7��|�i�#���@��v6Hk����7!U	��V.SN,�#ɛ�gsP�?�]���m����f�W���8���-�"(��π+���!��E�X���%~9V:!Q��h5��Ud�u%��Lc�\�5F�7@Y�'����j�A~��+�9���;r,2�(����6�.�@��-60�N疞�u�3 Fl��@�ج^u��]J�򑍥���]V/�,y�e!ѥ'����U�T�t��(�:��dٯ�q*C:�UӼ��w���e%]��}wZM���1j����{U�1�e��.?�XB�$* n���3a1���hoc%�S�.7SE���!k��t1ʬ�w�hO��_W&�NkI|��m��`(�S2:<%����CϹ:MʵB��~��̰�s���ze$~�Vr��?��������/U�j�������|�k���������As�>��i�������#N����c�3�H�{���ղ���|�x1��1�+-����qTzU��Z9�O�K!(j�IY~���sFo��*!%��q�
$B0Vǟ^���˄y[�]����z��c��幡nz���1p��r�^C^��ׇ}���	�|U�F]n�,�P:"���2���#[�؞KLf��1>�zRI)�S�}`����X	�h�4�e��+�{%��|K��a�lQ�[��Q����oQ&d9��ǖ���c����&��\�.7�C���>)ָCCry��K���u�<��c?^Wy+��&�-�a��)������J̷Lz���}h�|�F/Tݙ�O,���~vA⨦Բ��2N������H5Ġ�dǀ� XlE�O�w�aޮ�OV���8��>X�M�z/ٞD���#��ȸL6�z��D�}H48j�k-UŊwId!���  ɤ�W�M����K�׃{��a���.��.]Bi��`"�2�_����'Ar`q�����>�E�ԋ��cx��(t�8(%��Zd�9�J�u|�	ԇH��)�x�[QL,]ǎ�w��P�'>��1S1y �D����6f�Ş����}�ק��vW�\cޣ� ��!��3Rr�h��h'��|��o��I	1;�v����,]�9�E�F��f��U;�	��N�dN؅k1⥃K�nU���rS#�`(����9����咆zŶä8𣩏���/�}������B휊��ɝ[�3E$I���B�����霂�o²�P'��%�zf�����d�cy�������άUPYA�Ocfy�@�Q ��a�3�~�໡?gY�d�M9qa�WY�/ݢށ�1o��&x>R���������y�O��`�I��~��d�%:�<���Ɓӗ*v���M�s�eZ��FX��5>��✳֜,����%���S���9Op��ڏR�E�-���������@:����F�����~��%���b&�[-�v� 螖���q�S�{��ץC�V��h�8�n���p����g@C�u!"obaG`.�%���|��0�>��'n�)�@��/U�-n��-v!	�A��7lѿ��L,�K��!�����H�B����I����P:�?�GZ.}r<j�R� �]˸�����'Ư0����1��i�)-�Ui�z<Mr )b/��c` +\���\��|G�Շ��mz�k�t1w�0hl�ɽP�s{.L��b�\�����ڭjo�J+�_&�/�]lI�.t�]1�f���-���1qG������߱;�����Q��m/Mv'�C�4�vU�ݐ�������gV�~�jI,bw|��0CL�:8�aq�Ǐ͠:��bf����T�%���=��ip7�ԯOم��X����3	w�i^k{9��N�I�1���Vns'u}2[9������eⒾ��YF�GZ��<8-C�Z�Z
��q��˼��\��,��udǎ6rY�8q�����[��R����,Ka5E[]��E�e
��҄`��Q=(�/9`C�� ;���.�E{9�������A��*u�u�E3,�U�µ��h��R0?1����gE���^�c D��U��P��=ͦm��϶��n��!��?LAbX�8}��+v�*��'TK;���falScg�r���򴈺O������d~AW��3�����*�W렗�b&d��V�Cd��WҒ8?
;�Z&(jx#�JMj��d[�<˃ߡ�=\�]�y�^�~ŢE���h��^�F��Ł�����4"�$ǲk�4*��H���9�-%�ç�/��W5�����fZ"`e�
7.p����ҢJL��uf3�վ�,���;d��dDc���L���E�~5��J�R_�ƻP*{��i�K�N(�4R�a?��Ό�Z���I|��[h�X���7�E���3�B���l��a�8�-uW$&齯���1�����o�3��k��8@�Q�y��X7��ha!S�1q-?M�*+�3��K��X�-�U����xD�3@>߸/e��Y�Z��!��"��ew5Wȶ�f�!�Faa�K� �o]ai�;J�}ME�U���$���#T�)j��@s~��å�U��&�W;��Ҡ��;��:�=�pE�� 5� �0#��V����k��.ݦʲ�[���sR���1T4]�wFg�0B�o39�Q��p��ӳ�d]Wa���<ʮ
�C̍{�Q�g_.� �n;u��Cw�����"���InA�x�����ǉ�����!e��.M,ղ����5p=%B�%�-B|�0)�������Fa�j���I�������XJ�9���3��\<�{���Ef�Ӄ�/T����
�΀R�;��d�A��x�_Y7�&:��߲�!�cjv���T�\�  3��n�r����U�� �&�ذ{I�I|����[!Xמ��k/%��W����۟�GȺ�����n�<�b��g>O�5Z���v�PX��	�r<J���6铞�͢Wg��4��dw��>۳���fT�-�Q����+Nz�>Gq;D�O���rꡯ���e�7\����Q=,�Z�z^��p>0-�ߘ�#LXд#@��*��t�0�����@ \B's��2��օf�[�2����Rg%��'H��Y|�Ѐ�`���"{QlH���2��/�\�n��b�qZ��ϋ��#�R��V[~�F_��u�[���u7����a�Ӵ�Tx�#RM����6�gD7u���爲��t�nn�� ��=�l�}�����3H\���V�Fd��������ҝ� }HXm��1���Iª2��@jك������ܯ*N�0?�d�$���N(a��%L*����1g+3��c��y�R�k�@v��tO�%����ΔIp",��o�hd#�XwqTy+n@��u�1�x�>�a��|�ڭ�#1���X�v��/C_SZ[{|���FEv2��Wj�8�l�C�_rL$�L�Ry4=�����b0~����ԀZ'�*��R�ޔ�,^ݽ��Urc� �+��;������`���K�Xn�w�i.�_���y��QT)������2����ڹ��0c�U�*k��	�`�˯a��َ��vA>Q��GM�:}�Z�J&�~a����/g|9e�Q�aN :�Ǖ�&,2h�B����`P�X﮵����kdW���)8�p��X㙱���>�"� �F!����x���J��i�V�[_ZsW@,�=j����%�ۗ��ݍk����ʇ}�LbѼ8�q���g���W����]ڀƲ��2JG��	��e���;���A/����`��F��\���jY��"_~�i4�8��<�����V�����2�ffQ�v
/�!����!Rw-��΀V.l��~��1ō�J��_|Q���cg_�=11���	;I1��&8�y;i�DH���W)�.}���?���ןL ��}3vv�д��L��#�F
��">$�D~�rbۈ�{�|����������T��1 Mv�Q��{��@��*���r����ke���uN'f������'(�zҗ���0�_Z�m�bx�/Z�n�����a�d6$ �y�M�U,=�gXό��wr��-�����?,VK������bA��!;Y�r3Tr��g����[�����X!�����L�k�ğ� ��ġ�@���Fс=P���~M/����Z���S���F�$�����='��,��"1�%�R~$Ae4��2s�z^`���r��V9�QG���l���7������Nq���K]-����c��EȳS%�X=>�˕��=�1q��*��h��;�"�2��8���DfO�"�J8����K{�N\)��PQ�����x��_�s#�F�.��{����J˳lbq�<��q���_��G[i�&ۼ,s��
���t���dIe�w������@��t^o9�V[oE'�q�q���u��o�k��$@	� R�r$�x���Y?T�[�q���T�����K��Ato{#�P�l�Y�xsuf���$6�7�)�M�>-�h��%���/�A��`������Y>l�����!��1���:�;��Uw�:����o�Mf�P��"�+�B�xM�WL?E1?��P.6����i�U�B�^�м�����߸]lxg�wYH��,^�� ���4*gf)R� ���9��z�I����5�C8��/��Y38H-F@o���2'C�y0������y^ϣU6s�.'w���{�oQ���w�f��M��=Ŭ]��υq�Q�����N�ו]aB {�,���R�[8�O�Iğ�&�>�����R	�ʣ�$��{3��~|5O2��+���c������t���v��r���g�.��'ZY�z�X��9�0r5-V ��<�[��º���_�[�	�'�_�;P9����_�Ŗ��Y�+�F���d4���B��Bק�"�+�CS�>�y�Z�]��Պ�I�:!�zn�5e���%��a�Y9-i�=�5�Y�']�<n�#p�6���.����릺F|kkt.�
�|'��Ͻ�k��6�ASO�tJf�d��<&ΰFp��&԰[��5��QnU-'cK&���ۦ/۳yH�����ay꒿iؔ�h����o�W�� Aeq�/$M�H5&��(򷚅!t��C�RmG�j�m �!�?�r��\�oq�q̒�#2�Ǌ����.�[�{1i��"=:-}�ە��俎��ځg��f_BJ|�m�x%F��|˸}��NE���xt��@�곧���l$Ώez�Ԯ��}�Oq�fK�^�ϒ�4��o����*��a��:w@BWw133<����z�ت�B�v\���.k�`�I�j�������o�U~��]�6B�r:\��klg�F���,N�s@�n�{V���[+ b������������D����Y�j���0� �A6���#7�5�y��}�U���2���E��Xp��Ʉ��6|��S$�f���v�׹=�{@H�H,Q�2x�PEԽ3���
�D=�z��iR���	Q����8��b�J��.;�%�Y��?��h��R���Ԋ8���r�)d[=W���w�R�����<�êy�*S�v>J�	�1�g�`H(|��4��g���Yx�	xL��ӥr��v�C5�������*R$�#�B�A�G�)B�&TW���(D�NހD��C��eH��	��v�e�Eq�U����
�rR/�W��0��L�w��gҿ][ϸ�rk'�Cq���3��y��ļm��LP��D�'�PɄ_��=Hz|���k�3NŶ��X��(I��u|<����'�E�8����&-�{m�ht���9l�<Iy��ݡT�>ۗ��Ǿ<�����{ƚ0|}��)�ĕ�wu)�7���ǻ�RaI�ûpy�V�@�fk��c��o�ϺY�X�|�q�E�'Y��^ll�.��b���q1�\l��X>�5Vx�~1�&2��S�w�S�D\S����]�TY�M"��`�#9[Yсm�j"��U��3���uJ+w���藀�*\lI8��~���edX� Bo6�Ҷ'{թa>���5�J9��&3�#C�X��-*"�w��bYH����U�BxC�Z| �>"ڹ�V�{m��h�J49Z��B���m�������a���]V��@Pp��xM�Sr�(zM����\����l�\o�"�(q�ˇە��y) 8�h^���]��,}k�V�'�~`���ϚE
)���rr�j��e>���[H�`�MX���ц�K)in��[���	�:`1;0�Y�֪c��}
�hM0��~^;BW��#QZS�h�Z{�4�*�}��Ӟa�44}oG�xz�eCs��"e��K�\@==7����w"~�J�pk�ȥXb�]ޡz�%��pP�z�P+��L.��G��>%'�G�КU�-R�# 4�b�Tɺ��s=�L����}C'n%��V�oCC���������BIoފ�b��9�_O�D;���և٘��a�]JxO޲~:��)�f5^�`*���BeK~碌�hH���:Gߵׇ6C��R��qF�.�Y&��,��[U�������^�`l+,:�K%�3�IF�N���r_�25^�D���!X��-xX�!x�M���pJ|�1�Հ�s��{4e��#�k��!���'��8�1a<�F}&���E���-�� 	߀�:��(����{�X�c����(]I�w�$=����� :B>{�@3�N��O�U g�
�U�̭�ɒ��(�!*��7ˌ�{6wȸ4�[k@�/�Pz��9��5`?�@a2� �J�B"dO'����	�ͨBa�x��$m	�0��h�C�������gk�
N������=ݮx�K�Iq�P��x�e@l7��
�7�S�y$�&���G]��Jj��*���)�.��+c!��9�d�ot��C�(�$�+�8�$�ȫ�]S��� ��[t������hB|�c�{xOH�
N�2�lyg��)�א߃EJk;|�l���?���E�����X%�Ǵ���p�� ��md�@�t����T��b.(�
���|���2b3q������P~TzS�%��L�G����#ʂ��k�-�O!���yN�;�1�D��� 	��ox��Z�v4t��6_� ����Ta0TG*y���V����K$��ͯ�r�pʃ��ſ���"C}�s����'� �q��c��&�����7��[1?/Ȝ�%���
�=����!�� ��2^�و�v�R�9Ѩ�-��21^g�˟�.�ju���x�͍���D�p��	A�w)�?!�|�G��trrr����$N(筇"N���6X�a8'ip�~g��b�yn'jL���t���ɚ��~Fs�9�_o����t��X7F0\˳@�ŋ�<|���_������ ����pe��k��*���\��փG���C��;aC�:C>]����S�y]F�����i$D~����:!ނ�-��������7:F/~���ޠ���?�a%�)N� ��B����3n;X��ސٮ�����V9p������ƹe��y=(Y�8�A4C��V�������5ǌ<GC�Ljn�HZ@�]_���uQ������f��B� R���~�h]=O��;`��ˏ��N���}�Z�"��5Y��6�]y
�V6~�T1AҐE���%M�hi >���C�	eX\T�J�c�)KѨRM�����0�R��)�i3����!%�Р-R�v�y+���|!�����# �l[!.jV]��E���Nbhi�7)9��
Ƨ`c6y<ǳ�۠T���Ȗr��Hiӈ���k��J>��D���eñ�&7L*[�dtgZ�a^�8|鮓W��F����!e~�eO,|��,�H�$�̭�-���R�g9B�c��b�ݘ,��D�#f�d8S��>����d̄�sO^D�GIݡ�Əh$\hW��c�b�g�#�r="�N�������K�Ht��Kd\%��rV$�3^� ��$��`P����i�f�bh���)��C����K�+⏙�k1Bo��1�ZA��q�T����W��2˺U������R�0AewS�x@��Dӛщ���l�߲-�,G3�2�g�1�bgY[T
���u�T_������`�T� �eL�)���w�-��/z����G�mZ��퍫 �FJ>Ú�����4�� ^.E� (�I�e�U��R�I&ʯ�܆4(,�a6	�L��5l�n�<���̲QZ��%>������|i(�g�ӓE'�%�Ё�̼V�CaI��̈����Fx���ʷ��,�{�>�����)Yn�����o�pkچ"��E�e���/�l7�X n]%o��F� `n'�|9H��'�*��箼���6��!�(�@���CԾ圮���9�:�b�b�nǜ����9��VV�8�R:q)/	hc��ց������86:������H٭7������A�~q�@9LM���?�E���v��$�y���3N�y�z֋#8\������� �%¯�;(^(�?�/Gaz��Y=i�_HM�x��|'�!N�Y+�~�%E߳NU��������D�Z|�n'��r�܇5�V/����	l�~����(
%0�"㥲쯙.�'��H�� ��S>������g�D�vz���lW��-/�̅����ZL\f����ŋ�@ُ_sw7f�.�hB�#�#�BC5wiZ+�):ȱ_���ayvHQ��X�\����m'KF(J�ψ�vI���j���e_�!���9I��o_0�TӁ	�x<D����=4-�)�;j������S&&�S6)&����!9^��zz��J(���T������;F#[����\��q����@4'����r����m�����"NYwP+�b�M ��?ĩx1�ҧ��Dٯ�g�D�l��?"��>g���a�3Uګo�8	��"b���e��/Q�rOD�s�h!��)�9T�� ����W4�x�(�eo_N_�bm��c}�T1�v����p�G-�����>/VO���b3sߕmS�0Y�\<(;A�k�KsU�w��r.�1��(�jbk0Y=~O��NP�v����vt+���NǐO�7a�b�;d�/9֒6��H�C}�	��xO�������7��!+��8?��o��N
��7&����
��ʒW矸��o�lu�,e���3uoX��!{+A�^c�y�}�+ �8���N���^_XI}l��a��N�P��t�f��l�֙�6�A��C/m%S�;�>�il&&�~g�ө�U�Ij;�����-3e�3�9� |'����fJ���-���S��4m^l�4�N|�#<����2�
q���9E�+�2onq. Eg�S�ER�<��;�Hf�4h�_���P<��5��)�t� �t������4�$�E�%4ȓ�kHv��"{�Χ��|�������R3m�F� u�J�/��V�ݟ����ǄFA~�&�Q�7�uqʠ��܄�L�ջ �
�hL;��R�$��>��>$�si��GP��o���-�Z�	��RzVp�9��'_�-퐉�3��'�f�Nn#�ad���B������â��-���FK HG���)��P$��]�N�Ş���B�UD�*`�xs��Mk��>3"u�;яu�����Ha�~o��'S���
��H�E�(/,�����C��ﹰ�_��\c���
���>���־�K���-Z�Ŗ�,�p���d-���d�ɷ�6�3r�su\D���'�|%�
 ,��c�H��(����_dR���������	2XT
��ۮ`��&#��ɜ�q]�!uE�]@+7�N�Ǐ��]��1,N5�J�c5Iݴ6����n	����ApY�C�au>B��y��"H!�-y>���&�}���i%�P��(H/窣 <��Pi��n�2��+��S�L헇]~�l�C��B���������ݜ|�����c,�62|�a��HK����� Lc�'�U�w��%�:tT�E%P��h�;�qQ�Ǘ߂�CV�W�=,���ņuQұ$st-���y���
ͤ�m�v��y�M+u�f�M�iq}��6%���8+n�N��>t����
X�p��v�,�w҂�e%��)�61 �Ce��C$��_��gKW0%v��9?4�r�Q�2�<�-���Kv�k�F���*<���w~B	/8���0'�R�n�=�X�7�R�y��~����s�ؘe����.ǳ��x��3����&�����UH�9��k{�!��rbN�_�1#|6Z�r����9��
}�K�S葅��)��B߻N�1���|���2�Ok�-Ӗ*?���15�zy���������[:���F0JhG>�eO~��zG�U����ʹ�j��M��u���ʼ�U�������lq>��䚮s:�v'���~шd�
�<q$�n�\���U7���u�F)D;[@��TH�U:��by�a^u-y$h64=��<-3@���������>;�Ʋa�{F��C;��09�4��Y��ǰ��S��~�"�=�a(� EX���n�B�b��>����货ƨO�@Ir0��@+�"�0����,X�L H{6���]"A�X��0���g=Ȥ�Uf�x,M�{�͑�i�,z�_{I$�/��v�=j3&U��pc�W�qS`f��{�]�áL����%�U�r����*��mr��:l$�vLo�n�i�r��EB��I/ u=���F)J4��]������y"���Vי��d��ܹ8���Ι`�ݛg���,<NSu�>�͝���RLխ����E���@�����*Wt��d&W��IQ�{�ߕ_��d�[��O�`B��C��"��<�¶}��~�Q��# n��j>\�~��PhS�~�m}�:^��AI�x�Mҗ>��J	��fb��gd��0	�}�Zo��u���;�]ک�=DE���7EUݰfF<M�QH���6��h��~�>#iD�e�fm��A���ՙ�XƆ�}��������=A�N9�ϝ��49X���5�޴v�šEe��9���p�zh�88� 8�sxB}�e?�P�&����	<;�o�]*�i�8��z��˳�A��n?	���4R
��q�U�#eQ#�d�����!9IF���$��]˰�&�����{�*uH}˿@�P�J[CZ��.u/��ޘ+h�E�� XѤQL��tu�}�!16p���t"{b~�9�����25TKVr�
A��֢W[�0p��a*��g���x����J%'v�{G뜧�wX�,��K`BA��6 ��,* ���n������ruKTC���6�nU$��l[9���s�����ߢ�O�����¼u_�Xǅ�Z���ɁuN��I�2�W� ���Zw�gL�⤘ȟ��a�z�Q�q5u�b��S7����061A���X�����Χ���f2�<4~������}�̼<2�+#²��	G�{d?0�,X�8j�
r�M�z�\Á����@�*	�8���:|a�&G��]���&1xu�m����_SFhHu�j8�'���q���K�^�D�N�����}|��惘�
��x��\�/V� �<�Eea�D5��󰫐�h"ÿ���Q�r7�ICV5���p���sHs�3y����@��H&�)�3�-<O�c.c.N������̪��>Q�n-}��	gV�́#��=�����'t���4oZ^(������/�!6�����f�{5�e ,�(��f���ʢ�&�|�n�
�ͨ���wDo�X�Q[��+�sz(=�`�{��S|fO���B!��?<�L�ȶ��@
t.%��5񜓭-�dj�j҈�2��-\sB%�L�'�J�q_X��B�;Y	�+�)��m8��d�T�q��yec������)�pܜۓ=�7H7̴Ŏf�C�x�A� �b7k�=�\8$�٨�F�*"��@#�H9Q�>�n�%�w\�':��W�Ǣ��k�NO�|�a/�O�j����M��*����A&������cݱ�/���u𬑹}#�������ѱ�d�))N�����\��Dd��"�w�	�� N��z����o�~U ��%�C��,6ݽg*�w ��օ��&Ӊ	`c�AD	J:�X��

�9H�2���x�M0�Wh� £�� ��2�?�6si��Naq��w���%��r�����fb�7��ܯD���
�j�)BG��W>�3���j������ةy�k���=��r4{�ت�[4��7.9�hs�X�F��ϿL���0n������mg����UqU�c�A4\f�*��Udk���q������	��%r,S�^�L��Ԏ��+�W�l큄ȗ�eN��	Ѷ>N�ȯ*G��ex�m�\h�abߪ��Q`��l�o��d����DGq�w�?���A�L�D��4�@�.Fi~Q&�ެ��\ME&)�c���r3��Z Ovr9��C?ɾ;� J޷�9؂[��mi$�b��X�� ȫU�J�z��2`7T]��D�9>�0jK������y4�V��ī�WOѺ�K�x�m��x�F�3�y(�
�˼J����!�Q�T��=�]�F��Xzi�(�HcG۹MA�֒!h3@
Mrߞ�bX��/Z� ���.:xqP���9��طj�����@#��
��^�$��#�Gw<��[)�Iw$���刪vsNT�T@l#M�� 0pк��� "�g��WZZT���=)�=?>��2C�l�e�+�x��4�
���o��	V���-C;#��� 	���aӡ;t����-w<07s�p�x��Q��x�~&��%�����1�3h��c�?g6�]<y$���V����j��B7�UP� B�c�y#1h>�5�� A�FpA{ކQ��ԑ��Ş����
�ZB�j�q|�¿�O9,�D|�����5�gZG�-X �q�3�)-�$b�p��B]`����*I��r�����.y�Xv��B����>���1���k�_ �:��9�EE��R��uzVTV*� ��
��WZ�� ��V�b�ƥ��(���/e�0_�nD�8��� ���v�-p�?p���<��|Y盈�(���tn�ؘx
�r���������X�ە`8�d�f��!�'8~E������[O5u���&����7]_9��I��5Vk	���젬��:6.jk&��oi�tk��#�#�[��W�_]Y��bPQ�� gA/��!0����������>1P���5�%���YA+<�KdD׉��j��i8��Rr��	�)��Wδ������jp����=	�'&���3&��i���L����-4w|��$ ܯ���4����UlbPQ���\K`̂iΨ�/�?�c���M�5����,���Vu�-�+���	�0�(�1z�"Nb/����B2����]���pȫ}۵꫄�\V|\x��z�&H̗̞�����}�5J=T��'w��J�ĕ�s߉����JH����������� ��%���1Z�F�U�C'R��S�	��>�:�o5���}�-~r|7�I����OA����s������J��O{g��.�<	H�Г[�5�^���W��M+�>6l4�Q�v"�tA��6�8��9o�V�e����7{D� ��Ɔܿ���I7�>�o�8�v�sU�*��-�k���_+aoj���8(3�XSG�ܚ��������h�gڍ��g��v������^���rYL
+��M���UdI *�51ݪ;(��I|��7��gB��c���PDJ09&ْi� ����m�����v6��bI2P�!ͼ`雞�p����:ﵺ���a�C�!տ���`Y6�`k���\"V��<t��o���K�,���g�l���ɑ���n���.j�o�;�N����wke?f�H�L���r'� 
��C���
��qċ�9mdb�2]9u��%BܪZ /�ӵ��IBZ�"��E����f	L��,m�@�B�4�PRA!8��c�U�|�z��� %K�U���Bו�sd���4��@K��C���v��e�I��%����E�g�����5����$� �%�Íe(��$�7?�B;Q��
���|�hm��o�SÌ0�� �B�F=�S��|����b��s�	��<�*�6im� �1���L$� �����P��|Z��̌b'�.��4��1q�l��<��h��8H����ꟆFq2���#LwV�L��ܞb4�X�
S5�G�'A}��a�d�(��C��B�"�� gD�^$� 4y5��Xv�|
�`�#ߦY�9L ���W9Kס�tT�E�������������t��e�}!�q�dG��[^K����i	?1c���3�b���n��	�ĳ�h�4��4I5���s���;���ljGc�����[dd���=��L��Y�z9f$�J��ؘ��P�r���?o� ��eXǇ�o�g(�<�c�,y�%]������<{�� ��ҥ���:I{�8���H���8_/�g�ͳ�/Z�eX�� O�P���n�Kz�uf[N�s�B��ZӠ������_���4���C��%;�ftxɳ�:��C�������p�+_�@���O{��A�16���� �N�l�d-�_)J%���e���`�JiBҵ� d�h"�AD��GF�a#8�#��m�6��"��rϠJ �8q}�5"�^1񋬠��OR��J��X$�ʾ�2ݧ1��;��3y(��T:Ơ�Ze|+�;�J��m��8xK p�����D�H�0?��70x�1�\�8i�*��D��=3�?˝������7�C]ȗ�bs���V�S,�T,qƌP˚;$�@�R�I�HY�ǾK�6zj_����ׂ��穨i���%E9��K�v�ʥj�a@���QjN��R"�1wƁr���}�dض�w�t��q�G�B���`�P�\�j��P%����H`�	FGT2+��ܹ9�-/T����(���r���4탨����U2�y�htSi����<B�j�=P{��^�=3}��UQ�cC����Gj<��b�U/�[��4��E�Jc���[)	�UԦ�����e`#�q8�/���';Y�ʩ��z#�͂��bs�x8�S��=.����E^�4A��?�/�@��C��K��	�heϖ�A�^�Yn�5B�*����Q��i��A6�Hl�I��,m;��XD�\�D[E�rrv�n�����n'-��C@$�7θ3j���Y���C���{���r��6B���ebAp����#�u!dHkC�1���7�75�x\
O����.�]�.i��O6�Ƕ?Jnh~�Y�փÖ\PD�4''�a�u0��8�_��2�-�P<�ɪh���.l
iy���||��=��1��+V�����A�@8���f4*Ж�H��|h��$�(Ae"0�p%��X��9�h������V~�R�,$=5Ɋ|�H�T��k�zN���`�����e�e�0M6�S�p�]�x���	�	4��#"C�L��X�ɓm$������8��>��W/�T"+B���$h�{M��zq���n��玖j�0�bt׎�>�7�	W���I��)T�a�6�͂Ti�=6�A%�)W̍ҤA�Q���C�P���>~5�[P$�r���ل��E" ͩ�z�/v넌_��2-K������"�1'#�¤"�1pѽ��o��GY���z��v�@t<m�>���y9H+��Lk�'�|�>}/Tb��.K�:`�׊����<0N�y�rS<7��v,'�9'_���[Y��O�{uy膂l"���-�M}W1��}3�,Rx|B�����aT�v\�蟜<�`ɷQE;���MepH����
Z08�^�&ݯ͠}��������$Kt ٖ]�W�i!R����>A�TF�:;dn\"xH��:5^��z"L	k������|XD� ��غ����:Q�˹��/젏-"I���pJc�D>�_Pb:Q/}}��ߘ�_�4����@}����)��0�����X�7�7N�֦<Ia��1�à�#_z�pTJܔq%�/��A��������%������a�Eƥ
�$�Zx��2���yL��u�����S���E/=��R/+u
�D��G*Dȵ����3A��ਤ^�<toG���}�Aq�e�\��æk��+F�LѿwV_TT��yf�'$1?�0o		�#���f��-~u�!�r�S�.|�V|n�7���U9ml�������0�
�_����:rϭ�O�G����>��,&i.�>pǻc�|��ء/���0k��ku�+�k�+N}P��ܵ�ٟ4��;�'���D
�(O�z-����:��-��&��w����Sp�/�Z�0*p`1Jm;���0�,��+Ź1��>/P�� {����K��Nv��c��M)S7��dF0��JE(��R3[�'27��<GN�o�'-�Le;�	���&�&���>����<x�ܟ��&�������!:�:�;"~� ��5�6@�Y�-�=pdR-}��?'��Ý�/L����R	�4n�aGs���������l�nh���Wd�te�,��_�F����	E��4VuҐ���(f�p�aɷ�s�2lLպA�t��N`@^йY�t9Z��$����j�3�)��C6T�I�(k�!UGa��fX�U�l���&U+ ��Z����5����f]�9�Eb��\��)}��n�?_y��-%h�8yM0мӆ�XsE1�0��X$���t}�� ?IG!+y�]���'���J��#I+<M�D�K/�Fq�m.x��C~rӀ��`t��\~�b��{���٧T��z�q���� � ���2��RF��Dt��8�C:Ic�?-�Fid��mP�O��[����eϵ���)P�ڤ��=y����/��d��*`ˑ* 4nA!U%��ūU�]��ʢ�/z�k7GJ�&�݌�URm�X�x6<0�����ߥ�N�
������H��)I��4��N(�\O�p�3D�q9U�AeK^)t�W�
�_�>T��9�9P����p%�7h+��noy(;�.�L!���!�Vw��*Tje傖��΍�1'+A�hl��,Q���"N���_�MӚ�����7���0��j �q��#�˨� �f[��C������z��UJa-�-Ҹ9��6���}���4�Ϝ!�a6-$X�QS�c f�֎4��P�S���i���]�lЖ=��֕�4�]��".#LO{Ԉ]�վ�+.��ؗ�y��v9FG�H�\�!n��D� (��B��u�X�G��3�D����]���< ��o�n�J��,�Yp9mD�藾H�7EV��X�\sj�z��<Q"ri���R�@T�P�W��gE �Q�)��c�p��#��lo�RP#��0����+9c<Jg{�԰D`YԞ��|�YD2_a��!���n��9��ˬ������H5��-B�C��{�z�>��{���f�S�,��-��d�ו!!z1\ճwL	�2��1��ـ�Ko+jv��^0���jKE��<#��WS�w�L��i�x[*����xg�YNF���'�yc�#�Z��豓f2�O���]�Vp�5����x�y�0�yH+�_��f��3�����Sm�v"=u�@�4S�T*��|��<�ͺ��q���m�~Y���(��	�ߚ��Ϻ���� �m��X��1�H�k��$��d�-PEAg�ɇ׸@�kd�i�C�gNL:��a�K��($x�U��Ej���j7�����L����oDjڨ�<��b����S��.B=7��]y��/P���E�_��G��	S=�9N��C��(k��5b��2Xz�Së9�p�i传+�t@@�8"�QZ��!�e�@��"����!�� ��!)����?*u�nR� ���!�y7Y N�r�����F�.Hp�ǲ�4j'	��K�d�Z�ǌ|١@c���)3��<�!G�7��]2}%V8��,���oBߛ3����"`�� �a2W������P�hu�&~3�b�qB�gBz��q�l(�H�q�V�^�~4�j����aG�ݒA�S��m�?m�lD�Q�X~2�&���tT3����&���E��eqG�z� �8�~�
J����C8�E癵�\�=��Tm��1-a�|q������j���-��F�:��-�2Oc�H3����	�3|�aF�6����`��L��>�q�O�?J��5�n  �������ُ�	E＜K�d�v�c<D'����|~ة��P�޿x߄7u'��](�P�6�݃� �q�)܇�͓�/y)�Ye*`�{�%��B�J"��d�7�W�hb�[NL���L}���$�?��ɳX��(�5�Y��x՘�3��*��OV��}(���PW��?������A1S]3*�F����G5Ma�ѫN�κ�6���T���~�@������}B�~�K\���:󺥴(�����8ƛQ��b.�����c�k$�c]j�]�'��S����t�L��<[�6�r�c�x��čL�3؄  U���N����Fv]]x&����� v�#{˸�?��ɍm��0�=��5��$'j5��&�� �s��:��U�?�> �<)Vt�@��Ɉ�#�+���}K�I^!��x��~�sc!L'?O�X/V&�+�AȌ��,~+�:�,���)�=��B���n�{k%b�9���#Z�$���*��݋�}�$Ҩ�u^�T�ȆrLk�~^�ҟ�����1m��lE�6
.�1��-ӕ��IZ��飸_�/��k��s4~_��>>�HM��xh�ʎ�l�֞ڒ�<-��l#��Q3z%�[|<�:��|"���~��hu-:��6�x�t~OO=�<V��|�CeHvi}�Z`A�5Ʀ��W�V!H7�@�(�N��w˾��_�]S��T��*Ԅ��NhF���	5
k������+�A��<mf�=�٥�s�&?����q�p�w�=u��ilKt��x#S2]H䤸F ���|�-��n��z���k"d��ٟx��s������m�H�|�0Vmb�|Ѹe��2�XZ[�N��wmf��Y���%b�#MTs�%����^��䄘sU�4CO��r%�~'��f	��p�������7�Qéxѡ�)[��E�S	j7ښ���ͨ��� 0�P��na�4�Z��L�.�!�edi=��y��J���i�� ��-V��]��c�����fc�Tx�O�x%����`��]MGY_�6�W+p�6� �;�L=:W��J�J��-���t�1�.���knXV!͌$���=����$}M��	,�k�?5��^�@�NK��v9�1�t}
�S�� ^U��`�G��r����cp�!%o)�H��h�`�v��fÃ�gũf��p��'��$�M�üu�.��<�U:EX�A���~�lL��u��F �Ƙ�Ž��8���7S�p�QE�r�7�>�Fn1$gSq��-+C�q��c�"�	¸�{Ņ��6�Ѹ]�ߚ�k�i\���j.u�����$y���3��;��qy�U��0
ئ���e�Ye��� \=j��94�?v�X�h޽�QI"�w7D�\(,���;xiM^�C3gH�Գ����1�|Iʺ�^���,.��P�{�����CJ4Y��<�H��]�T��`�r�yZ��{[��] ��M�ئZ����h#8� u� 茧Xq����/:�^�ˤe�y��G��<�˫���|T�ls�M*'������FO,K�<S�έ�	�G��!ۚ9�$;s�� ����v�)z�����!'�&�
ji�5��	RXc
Iu��i������5��m��V啻.E��{���S �&��:�p�7G9�\í�X2.�%�^Mq��g�4g��+�.˦O����K� et����+9n#�
����ANz�xUG�����<�È�����aLo�D��Z\y9ڗː:�0�=g�<m�j���5�B6�M�n@�j7��	����Ta�*��.�@���A�3[r~-a~ɛM]�$��O�cٙ���?p��.�!Ձ�_�r9w+��2���0�h�VU���ѵ�d�)Vm�΀�X�%va�U�U��t�G���q�C_kMf������W��<��O�9�3�b��Ф�v2�܋);[Y*@\��9�9#���p�(S���_y��iu9�W�Q%i���(�8R�i��i�Yo�e�K�r�#?w�u����LS2���8�����9V�[�X~/��J��x��>��\����<����w^�����p��k��s-"+�gh�2+]�u�����o�0�����TedA-jI�L_������V�i�0���Xެ�|XS]��h�T����,M6uJ��؁y��y$,M�� ����l����P=���U���}��3��J@r�j`d�o積�W�6��<�l�>�[� ���o�������H��4U�/�9]
���ɏk�|y�gW0� Ü�Nx�d�g�g<�f�Ϳ��Zttз#*Uh��p	��7�?��мv�������H�O�f�7���`�U�1Ⱦb�~�Q�u���u���{R�2�7����b!`>����úZ�ы|�������F�f_!/��Mb��̔f��?s���řGd��omPz�}rU�Op'E%�_��y���C�A.~���)����s�#��!��(���W�<�j�^�gm��'�Z�C�UJ�u����E��d>������-]�1k����̖W�@���Vi��F�lE�b�7��B@{�$��K��;k'����R;o�D��43
�]u�ˢ�0�`�&�������RB���G�\��"T�pb���~�"؅Ht��Î��� ?o�y���I��ª-��D�@�_V�qە�יr���^�<�)[�Y�i�m΀<�R
X��XG��g:�L�s��uxQ�����̻#՟ ���v��H������"�&/��;�����F�_��H��,�1O�R
�B�we�L�hx+�>%��l��X�.�5����C.p�m�|� ���>L�GmA�j���?&E��dO�^�t�$�w,V���썃%j�i����q������؅
���)[��;K��l	���?b��8[z��*�H����T+���$�)���!�	چ�r8�E0x_;��?e��(L㙣�X#�	�����s�ќm�������gR~�}����1��n�a5���j0}Oh|�L�~*� ����X�q��H!��[ �<�4�cd^+�qY�{�E�7m��o*9u(�#x��ߝq��};��G�{��d��a�.,X�UN�I��B 妀g�Vq<��-��d4c�G#�?ᮽ�M?+�:� v���_�!�KZ�`+���Z��+c��ஂ 
V�*�����ֻu��_��ƫ�-eZ,�ZU�,Xl4���?��\>��h#07����`��$�r�NY6&I�|Hx�8ʪ*0\��XG���R�c�؎r �T��C��H�u��T�_S#W�Z]N�Wj?l��>!�Bc�:�.S=ƼW�U�-0�2�<x2�f~%M.Ǚ5�	{�o���Tl9�t��k��Ճ���N��ٞ8��ch�7�׹s���ѣ��e���!W��̩Z�ʳ�t�̀��x���m|u$�Y��K$�o�g�zY��ݜ��8G˙��z���)�����/&[�E~��O*��m#�Z��A�m���~-��IdXB6��4��cԈI1_ۭR,�D��>��y����qjMPk�	���K&*��j���0},d�r��{@�6@sb��X�R�u�W ���L��������/KL+d�����4�5M��� <Q1�~^�$`��
��Ȭ,�ò�m�y7z͓[`��������֨�G��g��)=�� ��۫�R>���$��-�5*+����j7�l�o��h��y������"� �D���Q@
�2�j������Bu�2��G�f���c��*(��404�qy�i#��:e�����K��g�񪯾�>u��`'G�L��>cX/^)�r��~���V9�B�HLŤ�;�<��?t��;�.�H��>��g@(��t*�s�T�z���#�[jQc�۔�P��H�	M ����;}E�X{{�!&��>�J�`F��h�4-�9uea�nGC��N�\օ3l`o������<媹 �b_��H�f�|]�@7����!���J\yD�c�����,�@�ݭd�����f%����V�Z>x
9'��XV�h��	B+�W�W�u��^[���t�z��kF͸�9K"�� �o��)S��*� �f�%��U��ی.&���TG�����S<Jmr���lf(B���I������\G!���S����z�l�VH�b̄ߤ��i�	��^�;[���K22M���!�A^�Ļ���ɏ��]F�¡�@�����B&�R[u�:V���^�*�]FԬ@���
�}ZR��r��eKOT��5�5r�
�o�<Jsx��yyJ��Hv�-W�l���z��6, ,��_��$���	VbQժE�������΋0���ȶ�D���~���D��+��ۭ)Ob�7���U?�%��^�!�����w����a��9,I�d���3�IA;��K��U����<�`��%�L���d�7@��j ��Ɋ��Pc�3x���VCQ��:���1�\�n����d��Ի�����B��q�L����)����Q	���]�'����NX���Q�<�L^mOw��[C�]oy��t���B}�1�gNE�@�:��, ˔Q
j��k��fL�n�6�S[�����ڔ-=�r]qt"c[m��z�w5�W��s�#���P�^���䗞��غ ��XZ���f���8}��#��]�D(�6"��TN���y����R-�3m��O32 N�5S�{m�<c��^s��R?��(�j������@FrFrl�(~E�Jq`����$J[��L��i�fv��X��a��gQ�	�̝��R�-�J�QK��CQ���T�����hf1�O���,*iʢ�Q�м8�N�[�1�h<R�Àj_���&9��������&V�Ϧ�����W�9P�)�k^>��b�h��/�<)A�܌c%�x�Qq����IS;��6^��J��;�^֛�1e�z��V�KE��G�x��� w����I$�
��i���5�d[O]>;�[�(W�?�}N���ÿ��k6���Qy���H����"�����#w�w�*Gx��z́����DS|0_K��d+Fn�D��Xu��e��Hv�g�Z 0:h?�̙Z�~@�p8�+݆��Kk�S�^��)�*Oqb#���.%�8p���QA4�A��$�=Ο؊H��k[yo ���Wp���X*�ɴk?�3����Hmr*���Uߔ�(s�={�<x;�N|tq.03�r��p>�Z��M�`s4��{RHa���?�>���GCz��'�*�EUg�+���d��.[�E/�0�tߐ4�z�k�bI���}�+���5>����%��%���[v0�͒��ޔ�f�
������r�L�����V-zFRP&��[,���'�������7ug��|,�:I�7�fT�����ડ��`�R��F#|�o����(���pϹ�t�Vl���?a���Ԥ%�@M���z3����M����.�s��Q0Irꛐ�Q��K��HLSk�af�:v@#V74JX]/��A�[��!m�p�=�q��Z��*�����m���\����%��o#'׆%5�ό�.$Ioӵ ���LS�[��`�̧K� {���_"���S�p���e,O�I ��h9F��#�<mH��<N���_R�Q�"<����P����\z�����cg�����O�"Z���2�7�2R��\	9{(�}��[N�t\�A���)䧚�ت�~�:o����}{�6�\��g�.3o��E챭�lP	�s�!��%����끌G�si��'�-�an��q w�Y8��&�����Ni������0�3�Ƹ.�l�XY�j��%�I ���75��+�Q�����/)>�Ǟ������H�问X��m��*4��Eػ;Rp��A�_W�pT��z�Q(���)��Y��M������*�E�n�~֍�<��˳�P����J׫��X����{�"�RDa���ur��:�Sށ���:�g��WhF���U�����р` Ʌ��̞T�s��5��d�n8墰ϩ�fu������:ېy�Y��g��aa����w�������Ə7��Z��^�^�8�֯�la��PN�9�f�f��H%�|>p[j��}/����Ȩ1�q��uqRR�i��iFd�P�a	@H�VU�>��d��h��_�QEsQ����@�����Sj-?�����s6�f2���%n0�Z4�Pw�O���f�V=�&o�ޢ6�x9�s_n2�ϙ��u����г��6��
ۣŻ�S�E�!ӥ���G��f[��ˢ��[�kp�ڲ���;T4����X�|�'�X��
���!Ѫ�̍EA�ؑ��-y��4�hҰÅ�c�m�C���o��GQ���Gu�
}��&���{���?!���bG؝��8}���6|��������}���J¢#t�TQ�����/���}�D���2L�]H�n��蛷|i�1Nx=����r�ԍ�(��G�I� �^�8/1�[N���Ģ�_�uybg�G*:�*���FC;�O)��r����90��E�K�����5�0� kNy�#M��jْI��H���2������G�X��e'#^gקd�w����'��Ր�Ea���mE~�w���Z�Mw��I�ݬ~�
��u*�9���8Ԫ��
��/LIw�詍$�w��i��n��e��=x]��(��B�熡ޗK�H%4��T1e�&�*9��7���z���A�;�Ʒ96݃��s�_���ᅖ�2�f�|�lL.cn�m����}حr�`���'�vX�n�/^��&�T�݆G���WI���z%��|��B^���$Ld�/E�ZW`�iN��őE��t�A�����:��\�Zd��w|=��	��^�]�1��e�4�8����g�ʄ�_�F�h�#5Ӊs�ix���U,�Dt
��3ΚhpP4C�9&�n�n�H�9����^ӎ�v�'��Kx��Վ�zn��o1ڃ��G��6Z��|^z�UV���)V ���8�@5�yp?��+�4�1d��֠|+�rh��b9ӥ��1�`��G�t���x޹�5:C�תi�25��U�{!�Kz-�y���$��������	J��Qm!κ)H�
�N��|-�f��F=ϝ:RA������СE�b=|g1n����:1K��¬�9!���^��	�i�{l�`x�]��( q��M�ٓ����Bf�S<s4��{�®;�L9�f(@#�Ӵ���՚�.�����3���4?}�	q(���)��1�-������\���y�?r">£�j(�$p���a���*�7	]3K��Sl�f�𽌣���!s�H�Ș�Q�WZ�s�O��Bz�pocx����Fn�]�9�o=�scX"����l��]�/^��Kk�&b�i�#y?�"�&��Ц�H��	�M[����
�Dq�RR������Lmb�������������?T ּW��T�8�١AQK\�䛋��y�:V1y�P���4��E�����jYg�%�P�y�g6����`Z�O~SCRۛl�>B�����8��0��)�E������� /c��!�������3�N�Zb�u蠝z�ot1�e�V䑮)ʹ��Xj"g�����{����N?��g�����a�^Үt�b�4o�2V�Z<���G�bNo}�o%��{�A�2�e�a��8HᵯN�!I6��:8�I�1[��(��y��b�����hK=�0zL�)�#D)cڏ�	�Ơ�tx���.�6���ẹ�I�$S׵��r$F�]&��#a^����"{��4s���c,��+��JZ��n�^��֨_E�svb�s�5�溒)A��/���;��y^���@���P����C7�@9!�>r�VDQm�v������*@N	��4⨢c��U�1��I�n�ꮹ��D8gx�[ק!��XNŊ����q&���$.�e�S�zl��1����(���bn��,�,"@n\�X�~,��fZ}�G���;w�,���H~s�I����]���&��0Iֆ7�d`���������̪X��ç��r�	[�%&�z�a����'4�.+� �.Lr�
:�:��Hb�����[X���'UP|��MGQ�ެE$�����, 1�+�E%��óq�	��'�O�����}[o����n
pp0�=>��J\�K�m�8ʮ�>��Ew��d�UNNլ��i9G��B���H�I��]�[KJR(^xdb�+�@)�n�������V	����{�,��8�ˤ)%��c�J[�h{���`S?�����2���z�!�^DqKX���@��Ʊ}v�V{W\k%��zu��-�w�@6<XE�}_�f~ :����
'KYM �A%�3v�9�Ǟ�'W:r�6*��'M�^�$��(�.�ӅM�ϓn4�"J�ѕ�(_ک�0A.�n�kN�o¿o�M�4W��]6n#w�9>�&2�Ÿ�tDQ����x�����G�M*�$�����]��:�)V��b7��ͪq�dI���a���D�ߒ�np=E_��<}f��DZ.D_NB��X���G����?^��a��!�� ��k �%��&1���.Zb&o�y��\� W�[��3'a�mzD��]Υ����޳k�w�N�նI8�a]|AҜ���N�!�<��LM���FZ\�e���t|��0�wq9���U_|�(��qY�gN`�������VL'�拏�-;�`���!��"~GP!6����M�����鱂W>����G7��W>�K��h5��x h��-8j)Cj�R@����]�,)Q�=�t��o�(���z������5$)ǒ·�(ߩ������LUr�%���m�۷�u�0�#�m�*�F�W�=���8^�w����5dж�}/:�ǃ�b�2>/��V�%��ӤU�9���1����w��>9�W37��p���B1�+.Żh����	2f�36������\�mxi�!\~ [�����OEO(�Ϙ�VL���V��m-�:��m��|�ˣ!8�ݽ�(�j4o}/z�9QӁ�=ǥ�g��� �X0�f�=PcY�b��Cl����]ü���_R���mب��JC<)3�_ȷ�ވ���{���t���	����#�r���.��J�X��af��)�rMd+�7�,}� {�F�D�(]ĿC��!acJ�V�ƹ��QOo�ɶ�K�k�M�{�&��@����ʈ%$���T��9?`�u��m��+L��^�n�^���	4��mن�ׯA9�6HXz<r����,� �/�RN78��*�FeΉ{[6�ܴ���������U1�,��XA�bQ���3��o検��*-��&���Q8�%�߷�4qǯ��PF��0�xuXo�t��CO��G�'�ڮ� ������:6|O����1k��Ju}Y4i\��Б��$�ǻ�Ho��]���s��?�.�`_�ߠzcA)�Ρ[��5��V����	�Z�*E����o-Gh���ϲ�%�~J�!��Z�mODq�&���!ƈ@~�[0H�8���՘1&�H��F��z
�6��m���[�0v�r��@�|������"ڮ=�~T~{�ח�DlLP��!�1-M6|d �L�(�� Ah��~nz�q<د�+_=�������KP�Z΁efM�QL׸c��rf����:�W
&_��wߩC�OͿ�@71�T�"6�0�����n��3p~����C�?a�~�\WW��b�'��C��[6VkҒ� k�a���y�S�"��"Y%:��O�LP×T�(�j�w�����ߴR��V�H����A.���q3��˪�J��ː�<��pr��"�+�"S�`\֚H8Sj��)x��+z3gհ���Z�.��\=�,Rʹ>V���2.��q��r����*L4���8I�^f���#U߳A�M�ǜh�+�7K��*Dk������Lgؾ�.=�,�	�e����P��>�,�_mO��.��6�;�02�"M_�p��U`�F.�k]�3Y��xSô�Q8>�mb?ߓ�=�K�%�$�e2� Ppћ*�?��zO#q�ud���@=v/�|�>ĊN_\M��f�|��o�ŋ�oV�qu�%ȓC�<���obE���xTs���E��%*>�R�B��Og�7t�Wy%���o��f1;����N�ykM��� �<����ţB�{�SK͋�`9��J|�"�#�,��1S�n��/�7�<
W4�kX����>n�J��-�y������J�r��,�1fƕT7�?0�)!���"��YɃN���&t�#O{ѶRw?&v}��?������uP�p�s�\��fY����;��m��IA����J~�e�K�|���k��۹d����2n(�a{½Hn'���,QL��2B��{j����㌫�5�L-:�Ǌ��k�`,���mohnx�SӠ��5Tұ:��y��7%(p˙�<_٠��CV11���*��);U��a����a���M[U!}�ڗL%J�J��"Ă�Ft���]��.8x6N9��-XR<�m��� �)C5KY��K����X�tG܆��0�R8+ð�Q4�?1З\�z��qON�!G�x���d�Ov��.��P���C)��e�d!��` 4�7�ܝrs&�c�:����L��e�w�����䢡�`�"�/y��d�y��-��;#J���D�����-�Ҭ�
H�N�X�p]6 v�4����ɓ�b������ʲ%��ԉs���C1�8zE���Z�E����_�i�5K�~3�,�5�j�@�˵3�b�ަ� X�V�����,b�-Wd>�9I �|ڐH�c�t7p��.��-�`���&R�}�KQ����)�SЀ��.l����: :�[�L��,oe)��d�u�P�G
f `�1�kzF�Fy�~��.�K�.�^9}��N+}=wHR��ax�G��?����Pg�6��:��_S^le%r��lD��G�c1�R��ujG�_ɧ�I
��7>"�Qm�^�Śm��t�!e�`�f��3�d�+1�1������n�&�8:�I9����~��,.��5K҆"��C�}��:���Ԗ&gҜt��v�;ԯ��n{XuIw ��hu�i�O�@�A���txđ4ňFߜ�^�ӂ�.�Eh�����g�?��iX��Uu3h�`��D��Rǌ�t�̊z�͞��3Kn�f�U�)���a��:	��e�+܇iTۋܮxƞzFH�0�9R�345[�\[�hm"I@������^CFN������u��j�  6��9�_�K�a��u-C.#��%����{�Zʟ(O^$���L$�����*���>AC���nb�? �(=&C�����)x
����p�fy��tT�L�z��6\�Dn�&P���gؓ�eЮ�/��|[��W����1��>�7��t&��Z��"�Q`(�� ����3n�7����J�_޲��u���)�ʛ��Z��Ŀ���ܸ�@��An4��h�\ZK�7ԣ��Ns �RG��+���kʝl��)r2Qo�9we��(�h�Dzj�k�K�p"���1.�����^}�L킠�E���#걶U0A��U��0p��1`�C��w�8�М 7��x�8Ƶ��0���G>�9!޴5��2�G,(Q�K�e oE)燓�`�纻4���ܼ�.�Ε�Bĵ$c>^�~I�N��1�d��N�T�̾�h}Kz��q6��N��w�yCb����J��?NS;[�q7΅s9Y�T�D�q�%3d���!Fw�ޖR���f<�W\����Y�_]�����
D�Ga�mXJ�j�T�`@Y���<�A���$#�s:[[���x��r��籕��F�4I,��wE�z|���U��ҹ�4��&mW�{��'�����g.��2�H�h�
�2'��[��*IQ�T&jUT���~��//�W���2	Y(�aF�y`�4����M��O�[�(�<���g!
�����Di	����A{��;�0ךӫ��E�u^I�$�a��˘^��b}�&�_^���Q1j0tG1���#�)en�`�"Sǐ�ʅܬ;���R��s�[#�@���gac����:��
��ʝ�!_Z��>�ZM�hZ�;Xp-B�noЬ�Ģ5|S諴Tt�1��fYR��,����@Trr� �j/!�b�^�*Ԫ\�ʣPH������1I��T&�C#?m=�E��L3f7a:��X~�~�b$�V�T�JZ	��8V�4��G{U�| 	ݿh�����A9q��R�M�{��:�&;h�5њr���gt�Q�g`�7 �&9��j�`�b:xSJ���lw�QY��:,�U�k%�����m��������=xy��L��9o7K>��Q�b��$��®s
���*��@g`>^�S3��Ŵ����7������1�?Z��Q'�.}�h�=í���]�w?l�Ҧ�B��N>���p���A��|Cүx��c�8���`�2��|������d;',������:�`l{�3#z�1QR��%��2�괦+|��$*E���,p���5�FTq�t-�-�q� t'(��&��?�S������1"� ͍3��o74D��$:Z1�ԉ���z<0��G�DW��t72[qe���$�����+�0Pe�ego�sj�e�5pI?G��J�da�P�"��A�[��.G2�5ٯ#4o��=�E,,������jX�>�e�+��z[�f�u�^Gh�1��>K?wo�Z��{�)��BPe��0�i��.�f �=�^mq����?�<��W�޷�莨�K�1����:�����!{c�f�)ڑ�����V���K�,J���ߚZ�?�y��b�*%�^S����r�E���wh��<PJx1��GSJ�z|��|�E>;Ã�Z�XMg�d}.��`g��٤2I&�L�L���z.�$�Ka�(� �l�`&V�'��������U��xS�q�6�ĽQ͢�_���Lg�.��'İ����on�&�������T\����PQ.	,+�g��I��*FD)�w�B�&�cRV�a\a%�0N$ �Ftl����Iс�8V�{�t9�1^[ I��Uoݴ�B�� �8C����d�K��R�_3ռN��6��&���4b�C�ԝ�����ߗ��j~�vi~������b�;�k��EQ������"H5��sU�_0zN�G�������j�lTz2J�B��1�d�ysX�eG�[A��a��+Q)U�l���d̘е]�t+�<�+�JT	���xd(is���P��l>)��_���,`�t�kh]Tt�:��:�t��m�2�^��X�6�4G�Ar�G��NZ�|�����4g��J�$���#!y�k�zk�Ӯ���k��	7���2���UO�<�������nK����}�	�oH�ן��3�)ն0�K������b#ZD��r�g��WSJ�Z3ܩN�=��°�����u�g��f����ٰ��U.VA��x\P�����)juȈ�qv��X*��$N�<��������X�6؋��:c�-�����;�68��}�9��[=+�;���pQ�)C�xv��>(��$}Y^�^����������|FB3��n�k�C����l���bP�t�80ｾAL�.}W�֬��H����I.��.պ�PO-�ĳ�M>y��E���I5X��$�b?p��l}���%TGzg×��fǋ����	v	[e �=Wъ��gtUQr���P�!�+�.����¾V�k���YR.��t���ㅗ'm&rZ������
S5mL͏�45��������|4��PFv,�936
��f�p���X��ŞߢQ\;I>U	�/!υ���^�k�4�{V�Sn�=X�hw႗��9$ϹrRA挆ސ�_)�T1uQ�@'6��U	�hP=��y%�f�X��U�S�%K����.�.��>�r�І�P#��&�x�����l�����vR�,7G����������yI���]���6��G��o2�=�Ċ�o�\��@��h��v�p+��-̺��d$��.u8,E�R2Qy-�I8�n�pYKi��j�T@�{6�ֿ�w{_[�A�w�dT�[�g�1�6�'�о̲�_PE�;Q����C0>�6��er���,��w}��&�tE��_�/�O/���-ȫTǮ� DwJ
\;��"JfW��|�Q`7O_cmD�,AX7d��n���	6����
 q�0����Up�'��W=�/������>I��	�q����X[��*��V#����I�,.`߮dN^5�3�)%NS%�Lq�E�����c�ZҒ�ݏ��5�mt�����bIw�;���&�+��KY�=1y�MWw8�W @��"��7j�[�~�[��jl1q���(�-������o��k�ݚ#��F�4�&t_�à����3���8!�p�gX��H��G(z�ms_�۟y6&�q+��F�����WË
G
�3��eσcL�ۄ��=5`;����upqe"���?��]���{�Оd�@D90O��S��̓���b����B6�U@e��v��]w�=����Puk�z�9;]|��bg�.~ўN�K�R�e����U���GQC�S:(-�0�<��kGU�c(��R�d~h{��x`���]ζ�M��Ӱ@L4	�m*��#�L�h��,�S�u8&p< �T�Ja��7��M�L��0�� Hd����d ��尹�P�h�T�J�},�����#�q��V��@�8N�,�⨃�UO��䪻��uڕ�ˀK�Hy�hFHix���H>#kB� sL΢�qqy�:	�HEo>.��`' �(��{��bc���),:ˆ�wH���mB|���ty�.���fU]K�G� P��![�]�T��I?T�\G�����ϗ�k�KSl
�Q�xq�5�%
C���yCˤ�"�s%��(�h����%S�&�ͧ�E��4���M��%/�Ӵ�$ye� ��$p�r	���T�(�X���Q?�^�7�5�����=k��-�Ga�ĺ�D�H��$�����"�=�!���/���iB����8�����%�8s��P�=6�!t��s��	�E���C�p�'�5ť�K;S��{21�̡��v�oɏF��f��J��"������"sꮫ�H&�����Sn�����MW�7����_���������@Y>F�"٘NV�6A�+~G���j����֠!`����Se���
�Q���:D�l��4�~ԓ�}M�Qש�g�L�������/a�&U,���ל8e������������v���X�^4�Y40�g+���Jj ���[%N����V�b��p�n����Ud�����[%��.����	��J�lUɧ~����0���6��
B��O�	5�RZ���S_(���8�C �و����
�{|:���� � ��,[b�s�8@�Cl��]�ꛮ�r�y� �s�_�(ՈwB^��H�SE����sev$��ޜ�M{fἄ��^�:����mR���<�׊��,����F[u;�{W#�;<�@������ B��=\H�kl��H
�m��6�>���*+�S�OlT�煴.N���F�k���A6�^��nqˠIз9C�g+�����M(Ԏ��%�*S�Vf���ދ�_�	G�����3�tWnR��������F��*����-Ժ`:A��g��Wݛ@.|�q�z�}�GZS����w��A��~�l�~P����{30�Pۨ`n#�j;�!4�����b�Cz������L{q%cx�2\Ȝ���ΕA�'\�,��F� �E��U�R`[C�wE9u� X��!2J�Ҷ�M���t&�������R: ��̖���-�i�1W�[�ipHS�@�(3���PF��L�"��D�����qq��FO�b?�H*���z%���ՙ�V��N)�!
Ά��r��-�%�����]��y+||�%���;�i��rbܓuI/��V�3����b(f���E��E���u�����0������p(�J�Ӧ��Ͷ��I$�:�����g�a��B�?(������eÖC�8N�`æ�t����%h'�p>�_W̬	3��y��Z%'&|{&�B\��wvH�Q��/=��6>�-����N߅�,ʻt�c�%G���C�7�����'���h��݇(	��������&�.Fc�e��=./,�b�z��Ʀ=�NM��aK|F�[�Kt	&�)�#�x��߇.Ğ� ��U��u����Vd�T�������_�4��޶�g�����i�Nzts{��b�U��Á?�^����<VUE��&��^�{R/LlW/�E���%��$u��������z���6��P�5G�`2G՗l�<I �fmB���ˡ�<s��.Q�{&|�^�r��%O��bB����'���O`glq�[�x�Cӳ�u��M���4����/.(���=�~�Ɣ�1E�O����*�y�Ǝ������,aK���~����b��3k�χ ��������*�KS�� �]]	�/&&��v�|
A9����;�IG,X������i��_��{?���wӷ��<������^�rBC�^��aIg�0r�,l��!��s��B�u�}�m�\��p�\2oD����K%pT/�����V���I��1j��]�l!��L]n= Z�(S�{�tV�j.P�����	&Q|
kW�����	l�"�*,�,��$���>�z1-R�`ζ0�'Y5͸|����?t��9����"K0�n ��'1�)�k�1�q�ɑ�{�����PaNl�U�?�����O�`x�7��Y�3��X�CLo��_��W�pt����nj.�F�R�+l)�E��7}<��كO�5ț*�uf�&`��H���h`��D������Ԉ�=4 �����ģ�z�
�����m�����J"��F�����J��BK��C�N����T�u���21��e� ���G>=t��FR*�&���_�<���:��o��|۸� �G-�T�u�G��
JR�����?��q�����.w`Xc6����U
�l>-� "9���{Ȳ�����"�`U��P��l����\�?�35"� �Q��^<H��Ϭ%{H��]�.s�㬶?6@�+��)���e�����+p P^x��Wj�zu�7�{���!�m�N�t�d�-�wue0���bI���_�t��
&��p�XG��'p�wrʕ6�!��ɗE��=�[�~A"�:��K�Kb(4;�K'�M��D��A��JCEEf��^%���+�h�\"JYOy�"PMXΛ��ۡ��X�aH)J��M�� KH��²��������J")#ψ/�~�=h6o�vIpb9��~��=�o��>����C��(����E��ey��ӓW�q�wh�n�x�1�<I=�S��{	�xD=�r�������J�����ɱ�O���O�4_>^�zk��1r�.�	�.�ʪ��5��!�F�k�bR�F#���&8Յ�!�{-@�{V}�ۘ��}���e�����A��,����~���X�L�qkro4f�u��(�8Ά�_R��@��0���y�w���%�lV�������S�BޥE�1Y����r�|;�9�S��J���{�z��3h������:u������~^3I�u���و�3��[�����8�ʜ��ٳ��t�5������hoՒPϴ}_��z��N�k�@\yeK��@��^d��Ml�����l�U������?����ۚ�1֒y$n#��]gtڼ:-0�B��E5̝�Vd_���Z��0J�d��`8\w^���g\��Ӵ��s�%��#����?��{���j���Z9�?~>7������i�q>�TT�o�f�.��qTorH��۠7~�=#{6'�E��P�����f�$��B�VȷV����a$�2��9��֐�e�d7�26r=�mp��`���K�j�COd���J�:X���K��U��~����nA�	g����[b4#�(�Lӽx���L��L�H���%�;�(�Gz�C�4Ӄ�a�JU[�ҷWu^�~a�g�Z#�����_���LO�ZWB�ϣL[�~6��h���z:ǯ���?4��c�"�$&������D�k�,ln�L6g(L>�0n$�1�1�N�\�%N)ecx*��Ń��q��W���W`�I�հ�$_c��OV�K���bM�AϬK1(ߞm�sJH�����k�eu�K�E�x)f�W7>Ǘ ���}��f�uhx����p+��L����a�b��E^�9��J�ds!bŏ�O���v�eOA���3��J4;���m��p���킵�]��x_t�z&�;���,v���K��E������(�~�s��Jm��薸~�V�O�g�z��n�ϧ�5'*�"��l;4��A� �"�g#���ratx�G4P���汜����XX���-)6���2뿎��С�O�BP�}9d�d���O�̏bE�Ϙ�'�1fQ�4���*����)�p�N,������(B����h����=%
�ͩ���-�:�<�|d��Є��[M/���Fl�s�hXX�r�*wC\��	Vn�?T@��,�8�����^���?�pF�)����PBT�j����P��^B+�.~�YYG���S�����obM��ͷ+�¯���� �B<$�B#5	��3T��_�gF<�P���SO�
��'Z՗�sN(;�"V�J�9p_�����: ���P��5�J�g��c;�W�m�Y8ttl�lZX\%��I¼�=𿟭��9�)�pjȄ0\���f��Lt4�ݕ7�5R��
����<xNW����".���7�f5��xo����|i���mYzb�'�>��	���=�Q 4��dGɯu���=�_�	H�e.ѧP�$�#�m�� �����}J���Q4K`��ݮ87KLG2aZ/_{�~c5Гy&��[a�>b�{M?��=k%�;`@oC�G�#2o!}fin���	�+"�qoԇ�X�� ���³L0�������F�1�����ю�n_��=�[i:`�D���Z�(K���/�J��0\ړƌ���V処]1��(�7+������F�T0�s��H���"��D"���4��'�4Iϖ�IL�+1(�7NV�$��R]�`����Y��_�
�R��u.����I�8*A��f�LhVe��ڴ6@gi��f0X��k�S����C\��2����=��}���X��gi`���(�iы�2:%�1$�S%898�M��]�p���xP����5wŵ�}�}�O��}�-*L��
�_e��$h�v������r%��X�������*Ym����o��f�@�,�\X4�s"GjWh�f�jѝ��oHo�� ���&�<W�H#��	1�)s��X�U(c�m0�Ίx�Z��� �46��}6g�V�uOV]�E��%�D] X��ZW�j��~?���<	��_Q� ��<E�T��s�K]��T�?��9~s?m^&�C|%x0
eA{�~r���>BQ<��&f#AbB}�XfP��38_�7���)�
��r�$��o���y����wM�g���%5�d�k�x�2 ����ߪdR�0˵�1��7Q�~q{�!gᠾ�f���K�%���}���^M��4~Nzg1�R�Ë*��)������T|q���kwr�b���Q����O*�� ���kd�r���%&���p��{�S�@�)&���c�}��
*�6�%2�j�'^m�|ʧ��pL�"ݳ!��`>�<���H���=������PJ�A�	 �|[t��c�'��6���_ώi���f�1h�Q�vh�iL�7��eh�S����k��&�&�<}]�U �ol��Cda[��&�F#�bȞɤsu�Mb;����vș�b�x2�'��a���*���b�K�n��U��<��dgK��[Z�	{BsdW�Q�?@�D;Y��0n�-�dC��B) (1�Kh7#Q�X�G��7�r�Cے]�n�7�얒N�57����_o�]�f�CǪ����������v!磓^q)��X2�\Q_ꕞ�<�����jw�:ד�{wވ�lҹ* JR~Qx�2a�y�n���°��d �~Ӱ�.=�����P|zМ���W�4`������l�.��7�L�L�S(c��Oa�?T75�q������hM���4���}��W.�d����zf{���&x��IA����̪_#q1ւ���ʬ
�`�v���/c�<�,�=���b5��l�ms�b�,!/#M���y
:>;�5�ǩ"Q.�I�&+634r*zf��&B�#@FJ��ZL*�fW����|��!ۉ�B�,�06 �!�K��pr��p:�7�	o�V�~r�	.�g9�+�7%���P���. �L�Uz*�,����,3�0娟tG��է��|�/h1�e�e����0�Q�z�����8��s�c� ���y�w����>!���(&R�uT��p��k��Wl��j��*pA�0Ee���~�@i�gPQ�LK�c>�6 Z�N(q��l��+�_���� b#�YH��	jf*Vdx�vl	^#���?:��0��"�kR��0�+-��=onB�,
������pZ�M��\���4E��~z��v`������LZ��us9���rp�m�\��6oao�6P�SM�jI��K۰�P���|ar���W�����[����8���S�l�$l$~r��"�*ҭ�Eq�V�s�T�1�+1
DF; 0j�g-����[�V`�-�b,�&b&�a�1��-
�� ������JW�E����@�P4,R6�{�D��ԛW��\}����WP#E�ZK����q�ه�|zu����T���;,6.�����ɑ�����Oa�HܮţS3H� [��W��2���kި�@��0<3�\IĚ%�K�ؠ�h]���B�z�}{Q���U��I�<��{�<u��9�>��i@��^*�j���K�u��R�`q��ȑ�g�l�=��Q #��^��Hm��LT{����_0��
p�A�-��i�X�Y^t�q��F�qi<�E�˧�V},�C���ˌ�m������7J�@��#������M�g�]�huM|�tT��B2uf(��h<)ʩy�w����tnPY���(X��yƌ_U��n�M�@�rd!-M���f⵹���ř��u K��
��,��ھ��j{�6��C'�r��U?���b���>Z���N��ד?z ����Ajf�?8��hўvkm}kR�;���;�W6�]�˓=���Aia�=�~(8�z��ַ��K���p�%�6X#-Z�dh���w�ch���;�%�"�]Tˤ�δcSN�]�3^n�f�w������I>Fܰo�
��Bw�_Z���Q�
`�!4���h�V�ì���	*���MZq��mu�he��|-Q�m�c�\O��n��m�N4�YsФz��'-�����'��`�i�ș@\P܈��T��|�\L�f��(���b��fQ0�R����6-
a����cd�6�M\�)&�w~\�2�ß�r�-�+�$�I̆��$Q8�؃2?=M�� Ƃl�?`Է�\~��B!N�Ʒ��[�_FP<g2�v?]j>?4�A�������t�^@<��"�����s�Afj]�j�|G+��t��7fM]������;f�.�� ^�
$T�}�G"��)�jAj8�}���G;>U����t$�kpRCI��`I$�ǫ��-:�Ξ���c����O}*�*���b�o�NQ���<��*�u1�~ڍ�Fg8>I?Z,�??9bw�,8!w��"�DE�7�Y�ɰG��9*g�KcI2���c,К�y(�z��XhbB+0l~�Ί��嗭c�t�'�\���(�	�%�Y��>�{��e+��sߥ�='�l����[*F��a�aY	jv*���W�QUvڋ�P����9�����-��p�b�;�3U�_�={oc���t�/��l�S2��M]L��D��Q�(�|�� f��̅�!�(�d}N2�Dx����B>�xm?v\�vd�,]��8�x~�)L����>����OxO�+�
Ex�jy��`7XW� a���?9���j?=P����(-���D \�k��6�](��J���R9>�1�e���P�<	��	C9�>�9���p��gr]�� ���{����Ea�O��� &����e���aU�)��Y��S�ˤ�.���y��؛>m�^�zLg����Ԥ�/ϧ>6q� 7�"�r��wV���g$Rt{�^n�0�|��O��vo����}�R�b�^�xKه�,K&��q�K)�b�����4�A$K�Aw�7�dX5E�/6 %��/��4|Q '���3qBR�O���<:x��T�+��[���.)�e���f9�F�B�l�#D�h�l@��f�����ͽO��� �Ҕ�J�9�"ҪNKr<wc���j@��X)�$2�XE2�Jݗ������L3�|�7="y����I=1r��`�+�����=|F�$Cg� =3��B>��)y��|+"8��A�3�����È]�
�@X-��V����A�z�i��	#j�ȗ�0���	��)�����7Q\�A:�bc�ƌ;���ZW���&z9����}V�>�ty�W�($��Fb���B ֟s�S��s˝s2Y�P�~kr��uK�YE�j��QȎ�z��N��3���!��[
�JV}��FUo�������Xәٵ�ޝ��4�*+�O�*�!��f��&l5��%����0���&=P~=A���ݍB��oD@�6!���i�ñ�^bY4�I:�v��fS�u.np�^��X����k���3��w��������kh�>��|��$�!��-,44�UY���>d'�@��(��9SrE��Փe���c>�H,�����$�7�W��~h�n����S�Dr]Z�ge⚓�C+}!�S�4��߳@}��b\�:AD��C�]EOH�����=�d�Uy]t�SA���N��I��q�w(�@7&g�$���,hTx���G���}���b_"�r'��A] ���Z`H���ӡ���A��ӴB/�xJ���ÅӃ��п7��vW�p���>|몕�ҷ�+>���p�A�M��7�p���B�tS�+�W�Q/0E�]���K�
��q��h^� r���=\�[A��
��K��K���a0Y'!;0TOɔl�
^`v�nk�#��6(�j����٧�l���f翐�I��V-���H�;�B�k���7Sv��`��W2���� �0��{C��2y\������!��] D�1
q4���_�$���T�%�>9��vOݙ��ܰHX�5�4��=3`�C�\l��,[���Q��y5O�$L�5w-v���AYHv�z����˙�=��L��=q*���JPב��3�b��7�=����z�J:������s*�߰��%�`=�"E�ߟ�l�S��<�V�Chj�m~���r1���)�e_x獕� ��=�n�&������KV����+�t��$T�/���p+���{m%W���(�+�]_)!]�I�AC0A�O�w�\Q���u�u-j� ��:o�Q�
'��o��4�E��>U�BxT<}��۰��h�>�&�K���s�X��Ȩ��ʪ
�3�K�qD����7�5r_O-ʹz�BJ\Fd!u9!r�~y�93>������!u�6�Y$���eS��9�� E��R8`)��^~9�S?ˑ��������r�Sm��>5��EH-��a�t��Qs�u$�"r�5�6Q�y?S|r���$F�Fkӭ'��H����KO��/�A�z��#���>��H��?��ݘ��c)cDMQ� ��Qn�hq|�69���Kܻ
�6r�7?�5��B���*��������(�2Ԙ� ��5GFQ8m>5�`�̰)�Z,<T���j��6�ƺK��1��4������mH���$�Մ�`�gO�5�
���~*W��XV�zr~�ϹS�����o368�.����w��	�Cg���3}oh��:��?����#�6l��f�㛆V"ai)������F
p^z-����PYj$4q��k4pvp1�0>��v�Կ�rɫ���k��I­j��<��TH ��Lcjh݈���J:�ŗZb$����]�+�fv��8� �rL+$T�k8����i�|��㥨�1%3�H��t^�2���bK�<�F(�)�����@z	�Ù8�׋+#��q�qs��Wy����F6n�9�5����a�{[#���K�����␕Z�.07���*=#��)vXK��fI��U���"}g��>�$5�M�C[]�5�{}�k3��������tљ#3�$�*��`�@�+��^D�=��9�q(D��Y�NkKhYZxgT�p�� ���.�wZ6�?m	~p�ڸյ�Ǿ�h�%��@tQ��ǔ&���>�J��L�8�'Y��m��ҭ�N�$�H���Zw�f�+�0.�#x�ױG�)e�$c٩�v�j3����o&b^Z`s7fM��ň?�j��~��C�5ßs  �
�<H���ty��ʈ��oz[.���P�w���{�$�nE�\��q��rR�O_�'�m��Vy$��/&MPj�DAx:Q���g���n�i ���@��$��Yfo��A�!Oٕ4�cW��]Ue|�{�� �:·J��^Q��\3���PG�~]=6$a����;�u�P8}9�n�,@�/��?2���!�fAG��"ܺ�����m��T�Yi���d�j���VF��D��^��P�K�=��%�K��w����d1 f�m&��Xw�4��L��Pw7i�d���FO����渖sw��69�����Es-�D!��P�i��Ӑ��D*��)Mf���ǒ��.���'��g�S�k�3�Ѓ�W��SPT��vL����`�q4"�z��"l{����[4�����ֶ�^��gU���s�1�80�n�}�Ϛ��<�ea2��~ҿ��.Q$H�5��OX})@@<��FX�A�=���}xs�U�U�Ȟq����|������a4 �rOZb�-�Ϲl/oU�glĲQBJ�"�1nAQ�E�
6�t �|��#�����E�̳㪡�cACX*���+�u��j7�vN��"�`.O��AI(\N8aJ�=�=57�$��.��	����\���B�hF[�W�g��Z�"�6Ls���S,uC.W��d��tw�;���u��o�\2������7&KvEqjid$�˪]%3�l�S�9L�glI\4�Tge��jS�B�O�sB�S�Юՠ �KJ�����x�9�d��[袠=�{�U��}�Ǽ3pS@-���ȋ��Q�#>�����Ia�@�+���>�d�%tN�S� ?�o?+�@�k�{6��R)"��h�G�CC�U`��s�
R���P�1Ӯs�P�xV-$ a�Y�?���/3������}�Z�_���Q3��C��4d���	�~s1�1���8ȵ��K�o�A���m�qv-w9@�=j�%Ȉ���=/�����.��X�_)�w��`E�jP�6ƺ{���?SXx�QD��J͘/)���ˑg�8�KNd"b<<���>w�z�_;;a>��H��a�T��uԏ�Xt���n�(��>v�dbR����*P;j]vHso�&>u��Z#5p�d���a����0�C3��qqtW8���k�8�l�4��~�Qӳ��J�!�lQ͍Ƞ�F4�wJ�����m����n�Y l%KkRBh�q9@\�����@�*�.E<}���I`ȟ�k�7�0���a���-�F�������6�	tS&��ڰ���z�nZ��fƨ��Od}C��S ׀�A]��)�隲��#�Z����E&���+c
�t뀕Υ�C�Q#5���\5*�i^�΅�^�V�M$��!Z��?���x�(������:�v�1q�l��%�K}����%��\T����Q����#�Y���"W���j67V�Ҽ>R�7%
�f�*����[�)=t�>�+s�Q�;z�K:]���uj/�%|��#�S��&� �t�J�k�	�< �$T� m&5 e��)�0��\9ɨ��8�����It����# 1�4^P�J���������}Wl�&%�˱��뽾��w�T�����ڊ���8<(��=�0�frC��T`~�k�ŉ��:��ʟ�MN�O �'j�
 ���^bh�^߮���rh�U}�^m����8��=�}<�hdEo�����D���[H�g5���^iա�-"�W�1�V��v�Ӑ�q���zɖ�wz�)_{��3���N��`�8"���tV��(���FW��Um����'�0vMG涄��2���[ewh.�YU��W:�������x.��|��J�ǩ��cmiJ�0&� � :���~��>��մg_�~��P�oz�g�ofGl�]�^����V��X�{��)/�A�.Ey���l���U�>��� �MD�������M�������e�SB	6Mך�w�:��5��W)1����8���A	V2B�W�Yx�6`�TU��Ys�5lX�a��fD,�Zp��9�b,�d��(����6�X=�ar]�H\#�#U�Pq��s゙��#GL�n��[N�E�I[D���YO)<��1Y�]6\B��O36�s{`e({S(?l:no�X�G����}4ИF�ȰqD�u��enm���>�*�F��V�q���A���Q�Ѡ�jX�W��k��ZC�#��a�������3h=�J�&9H�/��c�;doI��&��T?��,ߜܜ�����C_b�S��_����U�;�Y�D�������9�����tlѨ
��ޣ����
`,������J�Ջ��D?��}�͞UUl%��sג`8���<!��iɩ���y ��T(��U�,��lSm�|.��ɹK�X��|ϮW�d7v��X���0��,�\W�
@4�n�m�z��Ԩ\;�+�w��l{"2�4��XZ8���� �N��=�ݭ��T���ػ.�̓ �EԜ����/���.q�U�M'�$�,�C,me�!gB��������hs�-�Y
'��������IJyfza�|��8���`�,��0�G#���eۮ���?Mt�N5q<��/QYʞ��┊�,��Y'�H�ڡ��xSBY
��OSk�\�eU{�"Z�^�/��mm�.M�]�בd)�y�`i��n���������O���z�Q�(�wm�W��J��*�F�?�(35��8/���A?� G̑g��R��#1�~�h���_x����h��y��>�P�j��ȶ|�&�������"%)~{�b�8�Uz��	�=���aa����|� 3x�o���K/s�RN_�_�8��i.��}h���%��ԔX=/7��z�\�DGls�#nF����������6�U(����;�Bd[2;}��������p�,�s�|� `��O���՘�c�����6�峴N�O�VB�
�R���]���|�$z��,�t�q��m�f崽6�<C�b�Z��|�����U��Ip�65�9W���̊��ƐX��Xԣ��Fi�AX��m�69@�������u177yS��k�k<���dVWk�o�4�{�F��jp34��� �5��靇i��J �����q��Ot$�Qi�q�^��o�N��/��r:-�s�UpÑ�+i��rB�����W#N�q��a�d�0Q��b��N?�<9��c��NR�K�AS<1���+6��Y0��z 'd�d�����B����;0�}% $�����]^N�Z=E�%)N�&n��K��M�Ѭ�rB~�N��]�m����!�9���>r͘CG�0v�6~�NIY�:��2b�)L�dBh����8\���,��mC�X �ȇ�ݑQ�����0�$JHH.��s����� ������9쑁"e(�ݧ��@�S�:���"����v' H�V�.��	�A�S�.�FxX8fXCx��6�F�A�J�&^���2��oE�"�O-!_�f^���M��:���8�}��� S$|��5)�m��~Q����-b�*���1�Nb4�����T܆��C�iLЫ�����.��u��D���M�dg���@�L'�u�Gz>P���5'o�@����C%� ��Q޷��F�p�V-- ��������g4Ƹ��4n
���5�Y�'dz�XS�̕�=1�������m~+��� �Huآ�<I�*=��� ^�D��L?T�ƜW�Z�Dƹ�vP������7?u�@��޺��c����4C��o
DI|�u�2��@q|9��E��i�x����!}��Ɋ�v��a�M���H3N0�d��kd0^��%�9_!����7����8�N+��V� ��]c�q�/�-��j0d��9
�=�	T	I������9������v�C���=w�<�C��]C�H�QP�����Na*��`	@�3�����)��^���	4�O��R�W���U$�`�(�&;�G��E4@�&�/�l3�+��~�:َ��ݢ#˦���ع'�������
F��O���:	��2C�E�%\���7/�5�����I_��㎏፻%�~w��
t<>18B�:yE�Hg5k�� +�b��Bx�A�||�DI*��p'-l��O�r�1J?Q����`=�r�����6
n��`]3\����9��3���6QI,s�#D�+d�%>�(S�7��v�2�	IGZd����FY����ir�O�C��r��៵AC ;�L�Z×��ލZ̏Bd��Xz��ՈD?��+
3���|W;6�̪�����6�9 �;O���7K��m�?.��ԥ6KJ������a���w��Oe "�%_0A�n%n�gWq�U����K&nD{�����Ҝ6#���o���ƥ���a��Ǐ��ڊ4��H$�-�o� l.bW�oB�|���B��<�Hx~>+,�l5����(�Ing����%W�*ô��i뒈Ćm\�%p��i;�*<��z���]G&?a"�D��b�+�GP\ϖ��7=1����1�Hs�@tg��T��.T��C�~.ȫ} >?��E^��~�	����C��jپRr��-e=:M�(\����Iǘ�U �_�q!�ag6��!qBF*}��N��ؐ�=�U'��X�����֢�)�9Ʃ��~OQ|�&�H���)4�W��C�v�H'�a" %nD"s$��Ȍ�-\�á	�*b��zrÆ)@D�#ۻB$7�pu����篠�N����֟^�:� �G��:ٯ��#Y�_�����������:�eʡ�l��"V�����72<Z|�� o�k ��⌞���yP�{���u��ڻMNP�6x����CA�7��ڐ���x�����	[���k�@�ˆ|OCCy�cT5�0=�	�h賘c�lLs,��0�W�������3*F)��F÷ҭ+��y�.j��Ҟ�|U|H�s����'�8��2�*�����ރ绰�C�\Ǎ�y�[߬߼/C�{�V$Vx�x��>�N�[R�6��\��jb_ �"4m�}�e���gX(�G`c��ι�Ǫ�M��v(DP^'�p�p�v����3̊[Y����/�w�d�| a���e��*��d�&�yiX�_b��8��u��mu�
GsRL����r���'�쇠�d-�̵;v��������1��Nd��:�n�?��Oq_�K��H,�X�{�o��x�H�&n���~��h3$�l�AtdŲ��v������u���U�9�T�Lpt��|�ɮi��ځe~�D�������4֍�u6Ӳ���!�����]��'�X�S��	8Fc��������U�R�G���F����rD�K3r�+�۴��s�R^��*k/;!�;�E�G��ysz�F�8� ���CQ��{Z��dTC�эnImGΨQ�Ah����~�+V"�RC8Y�'tAP�Ԡ���k����ó��~ӪN<uD"�Ei���`;EH/�$���Չ��u륕,��W&���|�4��Ɲ�`������~���@�Y;Þ!Rqr���l����G˸ݫ��%�
��)Gz��׈+�A�;�x�/�&K?��	Af�!:�t[��j�����o�a��֕J_sjx$Ef0=�cX	(��B��1Y 0�A�|ǲ��	w�&`�����ѯq�VN�x��%���P��)�?3^aeq��+!�s���6ӂ�ш�h�%�~��F�]��"�H"�o�� ����
�T|��vl�\2�/,�`��i�5lOP|Ͳ�啯c��4�'�^L���:�ɴ�h�.�?R�M�k[3<�P�4F}&���^�T�u�n���# 7y�D�����VϜ|$pLA<.u�[��^?��y���|'����0p�/����E���Y�y}s#�2����W~��8)Z�7���������^�8j{�.��(�Ɲ�P Pipa�읹po����� �dA�pK���t�7�:��m���4\�ͱ�G�p�=/�V|��u߿�`�zo����T̊j
�h���He������G<p���Ӹ�~1���C�=n^�O��gnǤ��7,�>��v�eg������ �J������]���e�C�_��><�T{E`���J�=d�=mD�]��j����B��l�"т�.)��ֱ
g$;\�C�8 �ZIS�c� �:��F�?����s�����bmRC^!���l�,>�����'�� �֑��{HP��h	�,�p�P�z ����bn��`j�ȏXa��y�ź(j���Š�D%[x���
Yw���x�=�.l�xYb.���7���j}1Us��X��/i? ڰi��H�k�b��f1�68�o��8<f@�pn�)co��B��d~�L^���I���0<�z�3����M����^Dی"췹!aU�/���Y��p���qDl����!�O��F��!\aN9yj�ڃ� w���*�}�+��̹�8��塀@כS$Ȟ� �6��{��y�=��T�ue;�x菛�������(Հ�G�<Уk����1*_p�V$���i(�
��!V�L`b���4p��y���Cu�q���R�f����h�y�?��Q)����>&�U1Lʵo�#�)�+>�_̌�LD�a����z���wY~��S��z�}u�VH'F׳R)V]W�\"p�b|X	ۆ��>��b�hq��utͭ��:A��a��s�[�,2j&���89 t#c�'�
��Ɍ�g���HI��a�F�֫��nGĆ�)'x
ǅ> �Zg1�vl��&�R��_ma���mϠi-�\�Jf�!���쾵3*6�}���)��y	/�B"I�:r��<���������)s�7�m�����P+��ǋˌ�V�J�6#6�v��س�I?�T��̖��-W�0V xOi�Pc���]���n�����U$��Wйj�5�������x�~���Jy�IXbڝJ�C+�F��4e�����RcmJ⁳7�I4����s/�+�����={%p�5ohn�����oF3ʅ��$����u�yݶq�5��(v܏?S��~�����9��4���a
z�����������9�:6}(�GsE����o��F�eIy ֱ��@� ��2����|��](ѿܡ��ۖ�o���}UJU��X��I��>�KKIK� �/8%@�PSx�:d�ZKu��+&�>���Q�
��W
s�n*[��nL�s�5�e?
�拗H��eШ"�)}��|>T���}�����o��*��P���Hi~W��jJ�|�Q�`Aɮ��,Ǣ�i�^�_���{v�iR�vW�!��/�}�MR��U	D��7�[�z)w�gq���/�������;�/[�Y�^����=L�s���s��!fńW/7Z2|����ӕ0TItƎ�n�ow�f��ڼ�tj�W{$��N�B�TS�^�h���Z�����@P�|�<ۺ��`�Ƌ�R_�O�R;�8hL�̺�/@�n���LJפ�m�l�G �!�E\�Cf���	���`��t��_9��<��Z1���1�Ȇ�Ǵ�
���Ik�D�k�����a�n���ʨ��{n���9)��W8���2:P�`L=U5�1"3�{�B_�M�l�����#��#��f��@j�O���vkgI�nY�6��g*�;p��i6[���nq���Dt�R��1R5Z�ҿ��*_ƸR�S솏E�Ȼ�?/dz�F�W��Jkǁh�vg��w6Jb�����?�γ�K5������6� ������)�A���zP����%/�b{�_�z����vح6h���㋊��vh�H�b_��/�à���P�
T�8��D���OQ8�˜�J˳��)����{�/"�̯���[�{1T��W{�E���e��CWW7Ev)2 	)�ǊݲC��^���wt����� ���4i�YpW�[!�芁Tl̗��5ZK��]�������y�ڜ��'(�@f���`�;!�qhDh�������Yp	c��V�v�Kޏ���G��Ã�d<]��S���c�R��r��nZ7�x8���Y��%�	l��ͻ�D�p�diD�Nm�2����L�9�����2jB�����rHb�� |�{�H�X<>07r4l����23{�E>����ԴR.x)<z��n�h$~ĳR�s�u���y_|1(k����Ɗ1�qŞY�@��pŵ��J���N��!�&v�נ�H��R�d��:O����|��v���iGۃ=p
IQ7;R]��V7d��� �3y��1����txc���G�O-��z[�������՗Gʿw�%��	�X�����f��`���ziP�@�4��<}���"�?���:�NX#�B�MV����{��#_h��̋�� ��S0O��<��`��Q}�L�f
�Xv���}��ff�?��*�x�C9L�]��yq$�߹����C=��;�C�c%,ј�����A�$r!P��!�@�>e�r�Pwj=`�9E�y����TV�d��)���Og}W�8��eŊ���h�r3�zRs4�/�4H��D�<升�:.�Ęud�z^*�o���l3��7u���x~8H� d�ˍ�<h�S�{� �&2�0��]�S"/����=Ԟqv�� Q�߰.ף�˨Z?�M�:���b�q��.�4 1.�B�i�c�fk:��i�jV��9�0 �BL�۴���r�����n�8]-%�����ɿg�Nd������%�l�4�>|\�E��P.�P��,<�?���a9����r�yu�Gj�Ϫ��Y�Q�s}1ry�2���I�B�ë�v|� Kh{���)��h�w���Dˬӈ�2'1��@���B�+��Ƨ�M6�'�wW����uDj�}�t�$�.s��c�ء��R��������P�S()�v����a��Z�ׄN�y4�J�B �Px�
/�s,����ژ�����&����mPdVy��H�,�-�h^��u�ܝ9��<�j~Q$?�iȫ�Q��"�oXoL*=Q�$����ؔs
�t?�*c>�R����T6~���>Z������bu��ߌ�ȈOۃ�ޗXn������N
�X�Y)�T��X������7�^aeI*8�<�IP�V�0ޞ+�{'�X?��-���͆#�w���?.6���iL��r5w*�� ��+��2'Nġ賞����Itg~��" ��y]���{���'wU4:g�C�39�Z� ��h��F���{5����'��8��Bة*��d ��S�k�u���T`�԰��д�($���t�+��B�]K���
	'��8�"�|��࡜��e�Y�{[Rv��V�-<�H4t�y��Wrn�*�ÙS�~pؾx�N�!Z�Vl�{�e�������i�5�HR��;�����T�i��C@4��d/�l7�<�,~��7T'pZ,ݺy���}��t�ܪ,Ь@ڽf��H���H������;�^;!D
y�]L�n6����w^8���g�V(����I����q9d�8�u���"���º��R�ң 9S.}.;Z�N�_0��o��Jo"�Zz���P��S�~��=�/�Ӱ��E)8�K�HZ��U;�N3�{n?*�'U��q#�.�*\�;��P�V�8��k��>`Cbe�Ա]�͒�4�/�r��&�@�0�ũ�5e�L+�(%��q���|gĊe.����Ӑ��-i{"��#�e�+��l�m�md
��u{���=�B���ћs2z���<���*����BЄB�򚏫�Zn�%�ñ{���'f��Wn��鯾D���"n+���J�EaXc�`�"�O'dB����a�\PrC�?�t��ȶ�a��*H���� ^�2`��h@��_KVqSM\o��ȿ��b90p��e����Ѳ=0��>ax�&��a�(�|��� R	�*�X.�\�F}<�A#�&�@or6���
�N��<��\i^^�];	(��_`�P�[�1��"E�)����V^�m�m48�(�����M�9	'���޷<˳h��)�$N	����0*	��ݴ�x0��E[��hᘷ1����C6j7#��GAx����\c�ΖB��[�M��D!(�b��M4:��U=�׍�e�Ht-�Iã&=A�:��Գ�J�����=�d#)����2�}���0oݮ��C����e���]���� �Էg����cu��6*��|zOc���:$%1����UH�r������qˮOE�G1�/�zo�Yaz^}�k��Aʊ{O]�D۱�E�l�o��f��-4�dF�N@W]������=��H�{�}#�ş3�s��x�b��rU
����]��D�e�]z$x59tj p)�+>-�A��1v���F���T���$,1�\FE$9?�x60��Jl��Q�T��B�\֌���f
�);����"]�G_Y��ƂvA�E���gc3�֗Iu��ZH4�ZGH~sK� x�au�H�n��D{0��̏#��FM� ���j�5�_�m�$�5����w}�<�)���R�L�If����l9�9{Z��l��Dn�T]l�a$v���A���/��1Lz�_���#I��&'�pk���$���y����l�qk�wm��У��?�Bq臚�#m��>�7q���_o����o�y�� ?Ck�Yo�g������/�1�|����b/(h��dӝ��4� �g�	����*<R<����n�y��D�j�ցW$_��꽞k������7����H��s�QGTl�]��W�����QZ�BB�@�[4�`C���n%E{����j��5�	��9�=֋^F���^��\�d�g8��D��4.�b���h�f	���!Y��U�o,�E�s����8���|0>���1v��(+U A��뵥:��@ 1^��)��
��!zr������L�\�y�w���R݆���7rش�-j��w�ůQCOUz�,J�Əg��\K"�G�<��O4C���?�^br���ڤ�<�I#���E�'`�C���m)�{�!�<_����i���Re!c����v4X=�y�g$�3Y��%|����_!�x��'!
xe5ם{��}kT�W	Y�zz���DZE��:��O65/��VSx�q�� �i���:��ZHŁ�YCӬPW�T��;�$��Zh�WYeX���Rֽ�|��g�I5�<F'�����ڈ�3�P��[����R�RyE���T ��!�b��Q��I#��N�����z�d{ ��B���_�����F����~B߻`XW�o������#)&1��4�N�E�'�@Ԣ��R���Xn����E���Α���X"�ӎ��GϳBC�&��\Nw��]9����JXq����6�i�0����kr�{�[�rb$�����.����9LR:R}�+h��@�G6-�T�%���<��O!��Ϊ�����L9�	/wN<�݇F�n��~\���ӭ�g/e?Q����\e�2���َd����O�σ�G)�$�7�Sv�P_*�����t��p�0a�rK5��F۳�#�� �����:�v�M�0�0cۥu�M�3�3������#�W���v��z[�#:tήL��ƅf�����r阩���������7x�BS�ѷ�0*J�؉A��j�l�ׂ�?��:�7��[?�aCW�#s�'�}I`�n�l@}��x}7']��yL��^I�jC�(:D%�t���Uofrh{�1%��ɳ�h�ŘŀJUI�0g�ë��I͠����Ȩl�Ȋ+��]t,�
ṛJ�6���6-�r��T%F̖�����<��H�_�<d��U�<��a,|A�:��!}���?���)�䘴3
��m�qv�.������S�|�E��5���0��k}D]q)����"�*��Yi�t<��]�KqS�u�=�yF�',wO��!�(��������s���{Z�L&�R�yH���˾�DA�M�Aw�&HmD��R����ZN{qU����b߿���� c����S�$�܍Z���Mb��{"g�m�,��lQ�$	ӿ��J��|\D��]�Y_-���I���ܑ?	�ǟ�-���G��?�e{�9C��O�S���q7?�x�
�/59y8�%G�ǡ^qO��lEK��i�F[���\'�e�ֲ���Ex�XB���d�&&M��ً��q"�W�v�SN-H 7�ݬ�5t����[��z���u�02�ݷb��k�)�Y���z"�k���*�ċR"%���u$d��ƾ�������ҏԵ���tv����� ��4���.n�-j�;b[�iJ4ʉ�	��Z�	��'`X	����z��"���[C�.qx#��~�<��#����m/t�w��$�50�9��4��凘&Q��H+�X��pt�c�b��Vhw���Ro��'ԹM��	S���b/"��FA��;'�z��|�Lʤ�¡MʑZ8�B�a�?&SBD$���=L��%ȀM�4Q9V�Cܴ���GY�8X�P6\q<��B� N
���=�Γ��[\H�@|m4(^'�{
�V|�t��ݦ�S��Y)%�F2��$�-��s%؎V����!� �W){���*F0�ځ��q����h�VӉ�h�P����z�R�5Q�n�Ӷ�X`�>/��e<��n��k1`?[�>��F�8%TFB'W�^ |	�Q��j��xA�D��Y���d�;fkO��	���|�O�E�w//`�(9(H�FMyc�g���1oNH��aqSO�S��B�`LЅN�"ѩ"KW��ϑU����+�xg��9}�p��6@Qʉ���(h���d��<�yZ�N��(gǀƘ�>Ze:�J��˃AN���>�c���ե�-Z|GX��2���{�Z��� c���b�#B���'KP]��3��5v�'���h�Bm�����b0��V���2�kG��K�F�
�!P�O�4VOM����]�=!�%]�r����q����c���G20r6Kni�\C��ǜ &�֬��z�K��W]���bQߣ���f\+����;��
ưLd�ԑǇ�>i`�ޚC6'z�3�z�e�4P����kj�- �I��>L���g���g��/�ї���E�8߽-���"��U޻��	ݖZ%]pw|�urs4�4�g��O7�z�ǝ�R�����[1҃���l�hBk�b�5�rǗ99Xr/���F|��qq��ae<Ue40�!¬�vIm����TNA��~��U�k���Tz���Y$��%�	�[��7n�M=[�'�5h���
�<�[&��j\M���.��I��GaO�E��e�y�?��������TcJw�< ^�$q����0ks'����4��|�� ��։KXsьv%�'T<�����/Y���(��˭�����֮���JY�sU��yU��o��E�(H�$��C��2:86��JZ�|��K��Ze����{�U<��&�)��.Q|d9�2H��$4�GN�c��W[<�8o�&]@�#nn�"kW��h	��X�0���0�A�
WߥN�«Ne�m�9� �1���sL�B�1,�V�'�+pb���%�d����Ut��Hӥ����v� $�	���F]i3�&{���1��c�X�n!J;m�VRbO�AYdt��9��4]�}�x
��	8K��"&:�*'�S�:��9�#�5��?�é������g��� g�|I��]q�T�	��A���,����%"����$�gSv$P��:�%3�2�݈��`xZ�)Ø+����k݇�=��1�Sj8^����hv"��M��8��ʚ� �n1��m�%�n�iת����8��W��l'NA�@w�����|&�i����r\�J����O�gܟ:ͱ��y��G#x��'��@b0��R��0ԅ*��aD��tH�۟I��j�݋\��/(�_5�jΒYS&�m���������H��+����i����J�������ȸ���k��"-�H)�j�a�9�W�i��0.���
�&2�ry����	�q�
��ί�Kd΁$�u9��G�r��۠���6�-������vt!�������=��$~o���HPmN��K�4)� �fYӈ@�Ps\�6�R~m�,�k؂��|1g��r1ɻ���`\�cd�H�)�|#��J?�m`o�Y���H*��s�ЙEs�h�Y�����:���������B͚?�bK/���;d�{;'�{a�^��`�`n�����8��=�oKd��'����mK��u�}y�8�5	�'�֙b��j�@���P)�;9���g04���gҶ�a�@y�Jb���!��7�y����Ȑh���t�3~]��Ͻ 8�[�K;ת�[ʰP��x�DW�~�Xz\Ӂ/Ƥ��Q;���OK_-��ӻ�ל]o����m�.s	 ��Q��L��K�����6Q�4r� ���(�̯"W��H�kq�?����Q.��%��ʡ�«�O�uZ�K�#�/�;"O��1�S���[�K��~�E�+�a�"���ŨV c��b{�P���TL�l�n�ZƬ*e]l��s�9�'B��;�սE��]�E;{YTK���fkx� �E!:�?���\1��2/؞�	C���5����t]�'�:�����V�m"��\w|��=�?�u�w^��n�!6M'�$��a|{HR�A�5.��:O��o��v *:���
*FO��X���W�Q�]�ݢ__�M�.{�*��GX���,�y��")M�S_*�b����"������!=��R�))�|3�T��o�g�r*�b�2�JORd�xԠ�NO��]�2��gّ��s�Sȑ�/Sf�V�3p��;̮�/1CV�y�W<�y8F���|vw(�̓��Q]p�[��� �߬ͼ�dM��
����5I����3��*Wb�re���sɲ0w �ݕE�4mM�d��w��d
���ah���V���֢��	:���م����&�?��*��H��(W�Rso�,�f�u�h��-!T���m�D��t$�B�%�JL���n���Йc��N�Y��]ʉ��kZR�$��؍^?�v/��-4')���L~ s� s�P�(r���g�J3����V�D��1��LcJ�<�x^����"G-C�x6)I�1�Ox�C7���[�w���[��%�xz�<(�$-[CA��)ۆe���ap�Mޗ����F���"�o�[g/�L�)q8�_9l���w���;>�9oV�*o�+~����|O�.��ɳ��Ό���Ċ���[�w����}, b���j��k?5�}`��!�m�����H��@8��"�Za�;R���G#\�\x�@^�;�Di`�B���ǜ��![~`t%�pf�W:%�~�=%���M��i�k���$�0�evv^��ǃ�(�ӂ���W���y�f���ŕ΍�2Eo	\y���Z����ُQ�H�Y���|ŕ}'�@e?7�n�W�����܊��|&ƹ�gV�����5����*�K�%�?XS����%9��bj�1k�l`�R���S%ȩeC��o�dq��K��^�����i��.{3����ǪC�h�ɔ��^��c�.�ؚ\�d��������)���k�
~�RSal��9��	���ڷ�)�
�ďv(�9zi9/�>	��T��&�����,QX����pI��m'n�a
%%0`�������2��7������ӄ�D(�<Q���J�����@첫��'dP5���i��z�\ҍ9>>T�|`@I�FPF�ſ�[��.�G!n��,dS\j�=B4�.�j\���n�1 .�/ �����je�L�ٍl��|ϟ�CZ�ac@�V[�3NA]�G�&W�l`�(~�y�K��?���С�ga�|�����1@�Uo�'���nW�GѴ�0��O��D��dC�Yܬ�v>Q��o�P(��G27�˟�1��q��:��ip�4
Q��I�Ҹ�`ǅ��f�"Q�s��h�*p�53	ѫ� =Ѷ��H5 b�v_�s���B)����}�hb[b#kY�F�LJ�a�1����?ў�_�O�<)�vW�I�"��1���k�b�M�
�^�l�X�ūbZ�����e��M���c9��Nَ[7���J@��5r1�M�������#�BY�f���V�c9�T�t��-�N=\�`�KO&E�B������~�?L�Zq��>��$mZ�G�B�N��<�{�'�r��˃.Y�G%?�>l$���4�T�$`D8+��H��y���V�5l��_-��f�C*�u����	���A�k?� �LP-�R�DT�{OJ���W|�U�
]�xG@�Z��� �Î�=�U�𛐮���_�`/�_�|}s�F������q,�&���u���%B�w��t�&��a��E��/1�ݧ��mc��"��߽:��\�aM`��x�en6�@,ݔ��H}�Lļ���ʧ��m�I�~�ѡ*���ś� �I��{�S����_���J���\����r���u'ڥ٥�]�R����&K!'�Z�9uJ�Et��z�J�DQ�LXT�4�A�o͒.}�!���\�?Y���ҽ�B�m��u[�������Ƭ��U�ܵ-���C{K�Zǈ�,�n�5�k�Z>(���/Jy*�uxSu�j��~��
���(rܮT���ĕ�~c�����,�I �:�O?�W��� ��0�\�Y��I��'>�"~��VefRt�7%m�k�kY7wZ2�;����ŭ0�zaD����@�&C(��������B$Kn�e�D�^X$m���M�}�Ţ���D�g����\
;��(�B��G��.EÁ����W�e����Z�	��x�F���}�T�H0B�)���C	qxŶ+��7K#�ANmA	ٞƁ�� �{Q�4�$T�e�t�P�Q�ܘ^U%�yl(�[9�k���H%.q[��?!&W�>þ�:ص��go�r�E?�<�o'��"��3��������N�\Ͻ��C��Nk�,vum�߯�m���f/��
1Jh�n�q�@���
�F�m�k0h�(K�K�^-+�y��{�/�yE��Q����7CL�&a'��ͬw̫M���hMkᡵ���y
�z�hC;},���K�;r�t�ʋ�2=�ޙ	��)��Xt�4�_Qa�8v�G���S�<Y�>�����mt�)7r_�ܦ+�黝*�����W�%�Z?1�ڊQ�ǩx���s�!������r�4\$�іN��wѢG._�<@X����ĉcbq5sQ�#"}��ٰ䝲�ʐ�ʬ5����Fo_���6���Z�e㒙'NBL�[=�g��Y���|q6;9,:����m�9PSI��%��8�r���bZ!����F�T�ݑ��7�$�7�(��O��?��fی�e�ɇŇZ«�G
�)��#����֞6z�c��� X��p�1*Wt|\��SK�S�������O�>jXa�m�Qm�0יd^u"���MwNW���Y�'.'9���tN�}w��'g��jun�א$��v	*��䒑8EY��K
�sE�n/ɣ<?���}>���[��L���y�ݝ�m:Iڅ��l5Ok��F(`����}�=�T��b�gq�Eb��ޝI�=)h�Of�;+�i��_K��Ps�B���S�/7��G*�J�ޑ�Ba�K�t��z���I$M=�hT�����W�q/K0<��P����	�7�^J��X�������a�����S��<�ܩ�]�:`��ɛ�r�s#��z����rp�a������������p�/h��-Or'�J�t	J�kH8l�:b����5w����O5�h��i,W5܏��&w��j�|�p�I�w��i�H���1"��>k�!�W=%Ѷ�� 1��I|�L��6}�X�ڤ	������_�7G-S�GQa|�㋫�1��>�V����S\�Ec?dOt�f}]�Xc�P�CA�o��X�s<�Mءc�<j<z��𧞠{�+�'A_�d%�țο��@��>â��tE@M��E��4�;N�E�a������~�9:uM��A�R��u�z���ɀ{�h	o�L0{>��Z�+�8=Iy�*>./��{���.2��E���_�/�q
b�[B)1�l��'D��� ��8��� ��@�~�|���S@�3I7��(Q�.TsF3�������0ʷ>W���P?�I~�7���wM�$yQ�ִ����G�O�b<�w�����>kl�x�Wa���~�8��=3^��6��]���ų�KJZ�"�<�o�Y:��*�L���èS�Z\��l�����������鯎B90�0��R�_��������-ܧ�<��dXG�g�b�{�)XB�8$l~<���ێ�?ЭW\�� &8Ō��w�9.�t�|�T�(��y�E6���J���-��-ǒ2�'q��}^�|{�������-\�ǵ4U�0D��s�LJ�榺>��n�g関��l5�[�<z�ܗ�-Z��S�,�F��[�'ּ����a�0��$	�{C��E��!am����\���^��o>0�"k@5�B�0I��k��4q��{�oY������US����tO�7-��d���IIP�4�5'�}�4L��Ƚ����tM#Zxae�6�>o:�z�U�
��Vb��p� ���mS�X����!>�X�<����	���YGO�����d���gn/
�ێ�k$��7cH��H�S�W��V�>'�jz�idM;G�#s}�v�1��86����)�7A���j�a�-]�Y~_X��� ����~�QfMSo ��]�#�fkO�K�'��4��+늕�o��#Gω��xrX�z��X�oNO��`(�6L�M�jM��%D�hdrF�G���k�vԔ):�#��/kڠ�9N̫<I&���<(��9'"�����譽k�V��a��~hЏsШ.H�t��}�[";%�����a��L��پ��f����Ǉ 7�|փ��1�骼K���;Q,<� �x[�e�}9�P�|/��Z�]�*s~
�W�?'�����,��*C{؂M� &G��n��XD�b�+��q&��Z�5F^�[�?��)�s�m����8GQ��2�����0s����( �İ�2�����zf�>K+VpZf�.���U_���?�1N6�9o�D�N:������I��H�E�� hI<�����$7z�SxTE���yf�wDm�S�ιew����y��Rfk�������i�&m�q�Y�ǝ���2eUFJ/��H 9��G2�K\�!6PN�S�_�2�{C��*�U=O�F��T&Οdk1aPD�j�أ/��'�@��r�}|�ط��{�^�p�Ќ�����d}r�����lrIu��IgyA���6E[x^F�M�Wd��wQX�Ut��npLm,�����z���H�c��>OԦs0�����Ҏޚ�3�79���6��:��N4���q_�mB�~˲Ԡ�RU6
��6>��QO0f���s�0?g�]_X���"�V6�}}J�k�b*Pո�v��OL���#����&����8J�q'1ɼ�T	�VU�^;bqMc�4�!��ʷR��V�f����bV�1c�1D�&Ŕ&.�����k!��ln�#M��U)�L�JC  �$�_~Iю)�z����o
�p�sLs2��t
k�v�NQxB���%Lg��!���Ұ�M��'�X��^��~謔�7ۼ��I11�J���w9��#DlI���<�>L���i�����%E8�q?5?D�/q{2h`_x2����Nr����/���z-�9`��Z���3������z\�m֒s��Ъ�@���F��Éi\�����x����q
�dW�1	���Ϻ�#/c}=z�pu�2U
T�c���nЗHu�pR���?=_A;�-��G�`�K������C^�e�����>���5��x	As�vʯ���#%2��ʡ �T�V0��7��U�qv �6K�(d�3��s���<e%��ޔpl�[`!�]o����VP#湓9w��!D-LNR�͉,ηV�>�'i�"]B� ��_�]��K|*3�'*������	��\A�_�tNB�w����{�@1�:�'i��qsݯ�ۅ����w@�y�S��^���#���D��Θq�홃�&���RC�e�&�̂�||�c�vfU),���j55]βٙzm`�_���ubڋjUQ������>R\���
jH��?��S�����L��53��q(�sc
j�3J�MBV��/v����c�C" �L_�2WI?����+t|a��XŲ������f��.��gE�vv�.��2Yi�g���������܀5Пs(�S�p�ov�e>�P5�A��o	+��c��>�Α~�ѬT�%����|e���1ۡe����M��!� �ن��HL6��Ay�(����6'�ovR*)�� w�),������3���+1�xA��.Ï��}�S�K>� �[�rj�B�t�~h.��G����}��P�![��Ց���u:J�.��X'ƭ��7���PZ����?$~9��u�u7���WW�Q��j� �7#now�|���^;J;$S,M+���v��j����-�.�wY~�pWh�c�=d3ҕ�%�{f��~����^R
���gq���#��j��l�{�7��դB��BK���빚3l��˭ӈ���ȯ��6�c{��/������ 'x�^�s�JΣ8�>��4*���sC�Ƴ���!�\�xl��jA��l�L74�(徤�tf1�&A.C�߱���8h$�U�\� �q��Fb6��f�3]�d�;������β�WMpߨ���&�@��p���m���G����7�K�U�bL��]�_�����1{�6��4�3	O�ꊘ�lD��@fg������|}��ڜ΋���s`�,��z@˴٠��s�j��L�߆��\@]���T��|n!k���[/��Ƒ˒K��H��s��ǧ�p#Ç�� �]��*4��rb��廂����u�{_ I��Ԇ$s#[�
�A����ͼ#�3@o�O��өzұF�҈i�u����i�π�)�\��H�R�z$ݱ�0+��󊖁d$���M�$v��"���BxO����&�3M�r���u���٪j��&{6�)x�6Qj�S���D�����(�p���c_���:�A������}�y����a��Qc�h�
�m�.ݻ'�;td����#	a����/Ąn��T#1�Y{�;�f]�1��%��ি��"��k�Qȍ�YI���^)�^�h+����Z����Cak��,@�f~��y�$�R	��W�Z��RI���̢�����`qmX~�;	Q1��xKN�?o��(3�� �.uExg�� Z���[���UI���� ��ϨOQ��SĈW.�	zzH�[�
w$�rt{Q%݄�؇�f�^u��0��,���dw�y��K�r����l��K�6�% b5l����B\��FR͝�F�,�L�*�O�������ĊT�ˬϒ���-�0��5|V.|���l`��s %N<<�N���`�.�>�蟿�<[]'2$4c��	��ɩA�	�k:/���R�ğ���n��p<y���������M�FW6�u�")V�O�|՝�2)˭TP�u�ԭDJj�~��6�7����i��V�v��C���m���(b΄�v=Fr�7��sEE���"2e�8XގE�6įA��&�Ա���4�3�Y[�V[6#V��*���=DFK53���S���ah2������Ϭ�D����Hy����~jY��/�K�G�W�Վ*�X��~dy���9��^�
�#W@(��4�.Hp�zU;cOS9N�,I�-p@dA�n��%��6%+�����gz��z��Y���Ft��"�i< �Vǻ&w���X�H�9'��\n���Cy���Ӟː�|�xq�d���v�a�,cز��(�*�?!���t��!n��'r��v��wXs��h͚x\R�J0+�?t�06��/��QR��t	�ם��+qh�83C�#��m
���Zy��.�*�c�@�ڕ�:�f� &%a�%�ƙ���fq�&(��۽`@z�8dϗ@J��j�SW4<R�v�5ң�C�eCӨ�q9�ӻ����L�罙�"�h��[S��M`�ߋš�A��
��'��a�.^�?3�]��N���Lo]H}t_[���>�O�8q�Ǆ���:�LaH������zW�X�y���F����������ו5N�&U-dA���0�f��L�u���|��7����d��'^��u>��P�觐Î������~e��h&=���|�E��<�U��W��L�iI8��j`�F�D�x"o>��Y�Q\Z��r���vp�Zl�m���,��^�uj�=�T^O�ρ?lݬg���y���W̞�� 2z߻�0?�>�C���$��1�X����!y���<*�s�|}#��]��Z�Q��P�!�c�K�o��'V���T�QM#97��J4i7�ʊ|_�R:�E�OI>g����Pj \]����S�*�\Ż�T�L�<���`}%g�
>}�)% p�^�~Z���ޟ��~�p��K����hg������l�	R*E�i�!x���W�1{�BT꫕A2�?�|<�xmj
����]��akx��d����q�7�|�|a�i�.�pa��kf��v^:]>.V����.l�< &W�J�W���+�dD�6�\82�U�'�Q.M�ϸknpr����������Tn(~<�w��U�SՂ�js�\*Z���]�wG������T�C�1�+�"B'*m<�f�[��p<�"���`u�x��"x��e���|v7��Z|��z�Z��K��W��E��'��ʹT�Bǽ���\u�N�C���	��M�T�tS��ـL����LՒk�}�>ީ�OӮ��:&����?�(�J<�z�<��K��c�pm@咿���� �u�(B��C�
^�h=�p��K�������u�@�-4���'�����0J��(s�Ҭ�f�78z��0|��3z9q�nlR�x*�֙kap9�N�r�v�&=�Q�\߳؇fQ�;wq��)!�|I��
�=UW���S��ե�њ C���$^���fB+:�!`
��zp��5U�C��L㌧�C�c��I�S��Q��
�ܡ���,>�@%�y�o�6I�Gs�w�\"9:�y��wg��.�uA��a]���y��ȝL
0P�<�-]v ����)^DM���6�	v���t:ڈ�L/=�[����� z������l��HS��A��<�?:�}���@4*5|F}-�<̐r�IKV��5�r7�u�TWN�V�U�":췳q�Y��a�s�m:Y%i^<��pz���n�f(O��m��A��$��{l��V��Z���K�,��oJ~K�Ƭts��ԖI�{�f��P+�r���W"H��hG�񱢁ꈱ�ri�}�TQ�y��_��d7m�	!���1�^�i'���ui�$�Dnu�d����p��G���A�<�,�}�� �5�D��2wWԡ�(�*�u���Ŭ���r����~p�%J���v�ܵNe�(oja?��J{�&V��wI�[N�;R��:K�GS�0]a�A��No�rWc���:�D�R��Hm���S��4�A��z��ΰ�v��~��IP��?���a�m�e��֣�2(7�G��C����z���kҕv�)�H|�F�:��8''���p��s1���o:O8^j��g�p��1i����	W��b�{� ���~�G��h���B/�xuŬ������O��Ma�� :߀�F�oq���L�4�f�bַ�Y68�`�@x,�՜j8Wε��ZY��?�3�D(��+�#��R�r� E�d���<�`mX�̑G��E)���{,���W1e���R�����WA��$����Շ��i'����)I*�np�R-���G�����Y�2U�l;)������Ku[��Ʊ���{�
�.�5g�@@Is甸�x�J.ⱳ=*��})�)y�$�y�tܧ+L��UjW=��~�0ѧV����
���E�	촾�y�|Y�9�ìw������j�Z��'���!��g}��ni<�ڍ�MX�v~mk��h������[n�������q�V��x">���F,���b�u~kB�����E?MI��<�zT2�A��R�,�o}�.�`�����N����{`|��1?���uV
D����ݤu�N�����Z\@�^o+����ɍ�@t�f6�5�O�⒌��Z��*\�a�~���5��sؼys���&�J42��ǁvB�fӎ��
��b��'�dS�掵 ���"�2w/A5c��v�I� �
}��o�٬79L�v}G@���#��`Ԛ�3I^Fz#����djy��(�y0�1��1�>�#�0�z�S�:%|œX:۱��Q�V&mY��>��\�V2�|��,�p�#8�,1z� O�m�5���n����<�R�䳝��zjg��P��Y�� �0�'J���u�� �l�}��m@�����䁗�ɱ���z7�}1�����'[�{��X]5�q'wV� u |����K�c��?��⤐�E�R{m؜�A{3[���Y�\LC�/�P��&�%r+��j��ǓO��}=<7l؂�9+)��ؤ��"�5��?&\�.�A�#\��������z�����H�<��Ȯ����/[d$F��	n$����Kƶ�b�q���-~ֱ�8p9O*Yq���c�=ƁQ���R�nn���P6A:�|���kh��onTw׼����q+G�"��[��i�/��=g�5S���F1l��Y��VDf��7)����BBڌ)�.�$����M�P�1�8���Ւ�m�u-�:�/�ɸ� �6>t�7�d����~�!��/��~�\��a�Y+�oXE7���+6�V�H��>�|���qu�rl<�fٽI���U��v�}�{��Q��a�%�>���>Ι��A�Q��9tE��-�nb���7.V�9{����e��Մ����V���~��M�4�g�0mB�� 5�۳m�Eo%4�����H�k�QБ���ӏ=PfԢ)|��G'K8 ���g4��Q�	3���n�1x�N������-��@�.A�<�`�|#t�3��+A;�xH���j�!f��i�.��@���;P�숚�����ˑv,bH�g���d����w����A����0���WZp�DQCY�~�v�l� �9�CE��bc)��ƨ%v�`�'�\�J�^�!F"<s���;�J�:I�a��i)o��.�2c��%�6�:����U����K$"U�P�}�Pʟ��)���m�e���O�m�T�H?_�����kh�ULr0��9�����0淚�#jP[_V ٝD\�����>�\I}��O�Vh��O�9+��{"�RTd��IP���`�Tr�Q���&)�G�G���X%�7��#�ռf�������Ҹ�W� �=�"A�>.��b�qi�RL���Ғ/5�̫<�xᩈaE�*�t�UC��N��ھ������E�y"�z�)+G��NE�����8V{J�)Nx�V*�/O����S��(�P���8�^�h8�!���?�t��	��Lؤ�+�e����o;t
���:!l�1��>籑�#�q��][Z��*���-�{�c�d,z�<G���((A�/~���G@�<��?�d}W��9�ZIH>7LmH R_40�Aeʙ�!-�?�)���3@'`>V�getJ�p�f�/+��d�V��X�8��2˙IcA��3�k����bx��4�M2�۹+�$��:$>��3�cmF۔�w\�{�		4nB	�dk�������<���ݩ,�h�$�3?R�?�ͤe��a;s̩�_'|��Z��G�d�\M�s��ݓ�i^ʳ���9����6��U��O�g ��)T
w����~���TÙ;��"?E�6�!�x�`���[�`�c�rO锰(��n��ЬO!���jBu�"�ܥ`l�o���<��g[ 
M!p��-��\~8�+�o��Z�i|:^o��Ȏ�<@�Vy���%�|�4Z������z�z��?�`�A��e��9;#���qq�Fc:H���9I�v��pj��l��%u����z穹�ԉ����O��@e�J��SC�밦@�uԥV������:̄ ��F!P�wK�=�������y�)�Yȉ��x�_�2����a�$�PX�n���U-��9Ԍ�ȉ���<|�8@�����F�LhΦ���5�����ZMS=�&5�7H��6i��O6+�b��֦��Y~����ׯ�����X�{Up�+j5��ީ�r��4�Zk\ѡ�Է�V|�B�~�G��h��l�e��g�O�uXٌ���:�f8��V(zo/D9�n���&����fh������I�0k�k���Φ�Ky�\����D�a�*]�R�����}�����[Q,��cPB�|e)cZ>�,�$Eo��fa�ҐG:(4���W�#r< .d-�1}t+^��6ȼ.Xj�O���5ʻ[Z5���n@M'���RA��|�m kI8����`=r�WC!Å1���Op$�; �(#��bc�N4La¹���^ns�n�Y3�7a�UKA��.��f����pȁ�Y�m������3es���eY�[ʽ��V>B���-�(���N��/2�|d}���x@�����M�Ъ���	Oeլ���ɻ�U�(�=Id&�i\��s�K� K����I>��GU@`�v�je��u�$�\)��v'�
�= ���vu+S�QM2JH3|�^5 �xP��@���e9<>��'Z6i��*H=cm%K��6���U�0�ȷ�.Q�U��1�1&�G�Z�4y�LQ�������.rF�k/%�m��ú��7��	�wm�Jd�����3RT���/j�Udl��^��@�Q:��%����y��6��̖ih�%I���6����ɻ9`҂ɥ,�Zm0Z��ΑZ�F:a9R����ޗ�(��p�]
��ou�ȸY��d�Qg�_��2��6egjڱ���3L��y���S1��H{ii�_HS�\�D�����O�6��枻�<s{�˩@��>����a��J��?!�,)8B�$�f;�Q�|���i��t���≍2}]�xWq8���/���v��[�6"�W,B�}���!h�<�Ѭ%ٗ�
�H}��K~�%Aݐ�[P��}+��m�Z�m/�st*�C��J$�g��a;�ƹ����Q��pb��紺_%Q���q>b��Ơv��D�%R����p@��B"����[5#v��^�_���n���b]�"_w=�����ǆ�\I௵�w��D���G��.H)E����ES�D��m��
؄��da`��ᆘ����@������Q�$����4!�.#`Um���X/�Ԧ�{M���� <Q�Uu����J�E����J\�,���B+Z�1�3��,���M0�	\�|�
���m������,'h6r���M���Qݜka蓮ySkH����uEhָQ�����ǡ���4cf����5���Տ�k�9�?�UA7��&����?�z���zAa���Ɉs[�d����8+�k=��9�e����7#ب�A���lW�����6���A��r������i��=�U*���saܴF8�V�K4�m�N��c<��7��Q�_%B���6�;5p;]ʆ����-#�y��	 �b�@���f�T�
��Qi�^ܧ��+�y��]g6�]d_j�?m�{���#�r4���ʢj�y��O�����Tł�3q������d5j9R�*0ŷ~��hH��b�n��J�u������ ����§�<S�x@�a����M�ݻ�w��\)ww�w�}��?j��Urg�c�zWI��B��.�=$�R�hFt�z�F�h�B�&h+D$�:���ֿ�NJ�Hm��������Z.<%�^�!�ء�K�$n�60f@�S2�ߒ��KW��#�����I��my��0�z,m��@�-k�\ߨ�h�18�+��n�u�H�6	�dŻ22�'|�״�$C{���T�����)$%���-�DA�fAuX�# �B� �#�� z�Y���@m�A	4�v��d�:O��b5�P�a��)��6U �W>�G�M��/N�ث�ZH��rN� 2��>��A7��E��ԫ>���̀QV��=5�D��޺�_��ͼ�����4��\�y��E6���Ue['�.�R9��5�w��
@�ŝB�0�!�X)�%@��s��<�U����t]�2�=�f3����2�)ވ��j�a������Q^�A��w�^�f����Xӵ��Mu�^�8�I-�1��j7��R�l�lH3 \�2@�^�r����mҦ�7���y`e�L�@�h�^���z��'>���:��=p�g�7���v��v���(a�A���X!�;�
��غ!nʉoZط�7t�m����;7�g�d�FY�F_�'��=@--��QC߭�u�G�ia=.�i��(]S�X�-����ݸ/�o��s˘Wϰ��u�$&0�[���6�7���� 2%0mשP�`y�d��u�Ʃ,��[��B'$���;���bG^���0b����=�*�],XL�.�\��f0�$�%9\�$Rj}��pk��@B<u�>����zH��/��\���e��HGTr�K�<�\�y%��>�DU��q�2�\�7՞u#�
��Ȩ^Y� u󔕇��'4|x�fN����C0����Z�`�)�����Rq�s�[�O��`��Tf<�O�XOQ�(��e6U��3����R/$5�����d�$7xf�g������(�~_�Q-n`�t�F�<��.!���"�|/����H7����-��F���AS$(,=9��~��f]r+�0� ����B��p{7%T[0o�D����>��p��G����sU0�$��?70F|����l�Y^di��	�,��*h�Z�,*ٷ���:��~EE$����f��E�>�i.z����1�,F �}��.i�F��R_~A0�ި%k'�wu��a�[��_�B�f���1N�ʑ_u%�o�gO�l2�饟���o^p�&���#��z�ㅻ�9/H�p>��1�t�o���7�g��t?��zz�$��L%�C=W�я��<�--��mԛ�����5P���`q�O�!=K[�Pߵ���@h¬�;V/����I�  c�-�0����%�Z~L�����5�"I�P�%��_=9��'IXǠ#m>�B�}ę����⯬0�0	�b �5%������50:�.=�p��1�E���k�)�1���a�=�q��i�y�Qc��+"�\_����	?�w����%xs!�:�G,��<�]%�+���3�2Ff��޾�)�@L�ėX�>�#�)ZK��W.�q���3�ȩF�dRĞT� 溳=�t����5�-���cmkKF|����w;DB4��Mt*�W�NM�U��\��"��#I�1F�B�@+KAJ��=.����)>�(��@�J���L��0�}���K�-�Ew��yź���y`��e���HhB�f�u�&"����Ƿ*�	� �(�E�o�X�tw���ð� ���:��UΓR:���a�,��^�4K%3���x���������z�9O��z^q`���������!�X��kz�t���������8S��S�%��y��gF�rO��������DP���G�>��%8�Q�$�8ds��\�&feL\�S�@�_����h�:�-��r��,�t��	&Ž�->�فNDuNOz�����oCeQ}gΥ����z�b�j>+{$rf�-,���J��m�(���_�Z�ù���+!!��((�B�Ă4H�]� ���ꋎ0��(��?�H��>��;�I�3{��@7� ��a��W0i.���%CT�,���|i�џ�<i^�劸Jc�-� ��R��
e>� ���I�H�C�`o���`��&� /�KڈL���r��k�����#Q��BPrzZo�)ِ=� W*М]\gF��b�]�5*�U|a�R���!�^5�pRk�«�p�
1�gi�ϳq��
���W��<��81��eCP�)%�͔P��롪�����( +�`���i�k��}V�%��/��n�蕺�a4�ݭ/��VeP�4sh�C#�>���I�m�uǻʃ����Vyy� �h�3��$��X~�w�
$L�/�8[�cD�e˔�U��fV�m�.ﯮI�e:����#��&�݁� Xِ�tO�u��A���L� ���%L)LO�U���p��x���d�q�t�+y��WN�؈�پp62��	x\�f���0�o3��$�ua��"h=,qc���{���ԝna����i�'��1�<�~W�{$��� [�篇�uKS]�
����\�������c+4���-|�L �8d�PO�vH���V$���%7
ն)��s����p���.����,��m~�ʱ��q�;a�f˱�����ig�V�?^X6&��n���Z;���RG4�s�J����>�Z�!�i~�����a��9_��I2�R����R�{�I��c����pO�]��lܯ��s-/��PJ���A��;N�:	�d���'[��U�xf�4��J{�l�\��5�N�`R}G�6	
��?�k�t'芄�xv}h[K��G�|���4,�G稇���֯��s�7�uؐ��Q	T�Q���z�	���~3�`p�p�������e��0��e�>t�!�/��M)�Q�#ȵt�z�~I�`�"�ϠT1MP��K#�01 {�)�)^`0���&��d�~�2��Oh�<�*�g�O#q�ު�9N��j0�:T�l������Y��]��O�݆)m���W�Brh�{���~���b��4�'���f���j[�FlM�!�o� �(���₄��㿰��d�t؜��#c����Y>\њ�(��y�z��_�˜�l�H;�.�%��n(e�wݐ�jّ�iJ�����.��E�ۧF3���\�/��lH٠C�LcY��T�~��)a Nڈ<��<��4d�R��t�<V����n�!�`%Ĩ;�<�>|Q���o��)� �t�0lL���}�_O��P{��M:��(�+���5�\���P�9�Uf$bF�����H$�F>Z���/��f��he��е[_)}��(J�D���3�Y���-Og�����Alm� �C����Đ�s 7����
�H�فA�Ŵkv����з���	���|6!єR�h�waNG��g�7 1;D_J�b�0�SZ7o>�wpH���8Px�2�u4c������,���O֩��JkT 1���P�d:��9�dc��5S�V̧���T	I�u���2��P�)ͩ-�;C W(��@�K�t�<&`R�k2x�A�����罤"��qfcso/���<�"��0����k��p���e��2���~\���1���<���#��Aͧ���b�Q�2z�O �6%�\�ƀ���ߛ����\2��O 1��	GW����k�%7O���֏`ۖ�]�0�5�H�d����N��J�����d���0�5���8�P�V�m���yM�.+q��1�Y�@���a�����)�4�V�}�M��F��,\]l��U�Rs���/�jב*���CE��/2�=M!�ǜ*�lGw��z�9��(<I�!vbck
d������2�߹�s�Z��MQ�g�]N�.z�k����O��6����x���8�����C[ɂ��0j�Z�6�s��Y�gx����H*�S��^`������f�ͧ����<!�[��������I��;S��� -�AG�&`%����%,�,��:�w���c�+S�?�K����\��k�|h~��t�^��b��&&a�����L=뙞��Ē�-`��K������~�Qfq<�o��"d�p�kAE���N����:]�G���>ՙj���3�cP����Zɐ�F|H���2k¬��c�5�S*o�ت�ӫ�eW��d���֜��O���
���h j}�%*x���O�N!��ͬOi�����h'��:���n�������<�b��}���:���;�F8��B���������-�N�Z?�WH'F�C*�h!V]��@#����`��5t
3��~����fn��l��+%�'���Fv}Kҽ�ʹ)�#��#��.�D����PI`��Jt���v!�S\��W��Y&�_ȹ��9�Ib43=��P�}M�nvM�)e����#c�ӱ&x~�34�5E���D0zc*�v���p{�� �/�S[�J��ǆ�w��LG��I+:����N�p	��b��rI��~���5!�k'��/d��/��kE�<��u��Z�d`+D'�6{���@��Y;n�鶪t�&��iiGR�g ��+nq���X�P���Nq}u��f)��C��0T	�s���j'd�*D�a/ǅ�\���W��n���QŃس_�����}�Ҩ?�T�;��sf܏VS*qX"�P@o�	A�"�QԄ��?�WM�;ǿo�I2v<C���Y�Y�Մ��|��3k�Я�����͕^�����9��+�\z��er����,w�1�[r�2�s�3���_���S>*N�2#��<�g�Ll�9 ��(�`uW���9��C[��]�V����>E>R9��������'�|y�,ż� �_����ǶP?\A���l)��j�3Rg�E6�<�b���9��!�RΕ(���WS�^]2�ި�C���L��N"OJf�Ű�|�I�~�xy���x�}m �D^<�z]���C�S�j����"�:|�[��q���͂Np��P��ظ�W*
�Q)������=�oCM}@3��^�6��F��n �oxabr��`3�/�Mf
g�w^R]dKʽ'H�U/3����e�`}�e�\�F�r׳<!�R;����"n�(:�-ӧW���~��~C�)&�)�Ͼ�2,G�Fذ����,�oh]M��c�/>z����9���Zzo�WH�O��X7�o��_O��Ϸ�?䬉ϗF�~��$��r~H�l�����=�3�L�cH�	
��_U����SA��f+�pt:��G�Gw�)�#\����^_L}���BB����+��j);�!}�_�8�ԉT}��@���Z���lB���#�
��T��0/���A�0Uv�U��Dx���k���DY��?�G�S�G��4hɢ��`.
N?�gXSy���n���@��W�s��I���gWSFϽ��������C8�t����	��z8��2��Y~rY$�mw���0i^���i��O���(�]����Z���N�g
�ԎR��:���\����*нd#Ͼ��!�>�s�^���uq���R�lG���G�i�[�|*Щ�^�Qg�T�
z�OAۄM���S.#�0���S��!���1�Q$�T� ��}��F��a�"�d��jw�C�_"�����	������,=��1��?�6�����U֩�[�ݾ.[���1�5w�,��y*}x����ɱ9=e�"��s�L��"���q�8��g�:���[u�w�o`(�HR�L�&���Սm�8��t�Z�Qb������5���	�	Ɓj����!zC��iÍ�����b�-[����1���=�j=x�}񫌒��"���QD�����uŢ���
�y#���F�:$��
	���G�fU4.�U|�b� ��f ��{I����}4����������9tg]]n�;�B�o.r�f� ����?�{�� %*0V��F�FVܧ5ύ� \���|��b���2�a+e���Iorb[��ѝ���M�)�I��u듲�,f}���[9D�$�4� �.q@�4�"^YY��J�`���/B!�.��h����6kyM}�5�nv����GmƛG4���A��0W��oS@K(۞���£�RT7�d��@e�8"���Ý?�xDq��L�"�?��;ҏ�`xˢ����>�� �RO���1��%�v��P*hP�Q������p�����\l�"oNG��~�d��v�&���h�@�\������	����6Q���yM�Jh���aۏ�����yZtD��46�K�LuxPyZ�.h�[���Sv���8��FoŜ��h,��H'�S�������(�������$e8o@l{d*ȸ�8�/Ɍ`+Lu  R�;|�MG�m ��Rs�29��
LC$$b���*k�9u]�_�u2�e���������Ú�Ἂ#�^���MBXg�����ʕ'z}��
�Qz-�A��g��Y
��� ����g�Mt}�-�ȟ=� +���=�6���6�h=�bGkC�aoӕŴ�!�h��<��̹W���CgBv���#v6G���	l�>W�T��<_</�X�{����S�qQ��
�5!�Q�e���O=6(J�,L�ʟc��u#����=#c[���P,�+��~{�Ŝ=�	�-�+��e�$�1k�fm���_�-n���\hJ7.�(�XG�,x��BԚs+�9�١����j,�2E��a�H��Sqvc[$�t�@y�3(n�=/
HM�P�~�$��G1�(I�N��_uz���	Q��Q��k���ᇖ`��"ҋ��'P�ϡ}b�rP�w��VoDB�G��2�7g��lvk�aL���!����Η|��S�����_p��E�cC��؇� ����,���焯1��A�Cv`;V�g�@K�0[�e]�6��!}K .�堏&J~���7H���w��ݙ���N���lh�ǂ:�/��^4?iA
��'~Ɉ�����Զf�̋��)�H
2�y?��b�t�n���2t0yU����_!����]"�6?�����#Z���}0��K�놠�+��X}XĜ���3��Z�V.�'�a�����,r6����-o� ����G�n�Q�l����+<��E������[L s���,��,ٗ��j~U���JW��')5{u�rM^�ެdP��v4W�<\�!}���x���e��b�4ͼ*�A�jj�)vF��wZ��h߆�=�,wv!S�
� �qx��@�ܬTM��dE�,�w�����cZ|5��:��k���3kS��t���*kFW��SF�-��i��ܹY��yi�>͸��qDS 5eoq}�q�+�3�OD����#V�RO@N��n�'�Jɭ!�۪ݓ�a�nN���n�#oW��KH�>/�!��_��"����V�;���t��nZl(k�#vr��u�X{e�d��Cb�vQ�^��κ�_mCf\i-H�)�R�x����.�3��e06RXV],�ؙy��Z����;��Ue��`���5�mrn@L� ��s�p�j
�P���<etl�b�l�M���OĿ�D����tе��O�P��CH�\�1f3g�R���_�Y��@��N�����L���tF�5��~r���fh
�x�d��C#V�G�6%E!6�T���LU�+��Z��ݼ���S�,X%��`�:7�r褰�B�B ��|zf��1nϝ�u޲:l�� c�Hgޛ�E��kIu�%�}R��S� C\�9G���f[���h[WB����<���6�;��Bq=���]l�����i�����ɵgk����u��	����,E����k�n>�C��.����xp�r��<��tP7 Yg*U���XR�}�D���Io�SV�ϱ���=��(Ӱ)��P��sx�w�uR�Ҥ�ӆ�3V�ABRBf��\�Ϛ�z1J�q�-" ً �|�7���C�`��Kd=��g�k�j��U����_���>�����o4��U7�Ĉ����/�s�!AA:����Tz ����ط��J �N��-��i���"��qZ�>��ֆ�X��sy��=b��-��'�G�Pȸ��c�ï@���ʸM�Mqkrg���d���=�"�dk��\����3l�x�&��w�P�o���z��>�&�I����f�C�I�X��$���1ܼ��C�ѠS�w��h���Vc#�O�`�u��m7rY�W��l��u򝉟�R�I����cr'-��-�����_�'�9*��b���miYt Xкu�H6@w�(.�QEXw�JЉ����S���N��Rn��J�|b]h�Y�p����bڕ���r����F���;��l��{뾠

��l�!��C��kʖ��j�h�Sw&���F��C ��n�#E�q������a'��YN�l�A�����j�rx{&�op�b2i5����z�B�JV�H2H�Ĵ�;�1m2u`�5��Z�r�Q�����=�=���D��8Y�0EL�Hj�7�jŘ����^�#7Z�;$	�'o�c�0κtr���r����X���g2K��Ž�կW�Gٓf��:�oi�&X��u �IY�:�I��uڣr׍��I��xQ�W}?�hG(l��k�_��<a���;r����e�
�+���I�]E61��@(��i4���/�����H��s�ʶX��6Ά��%��/�0��2p�V��|7t��R��ӑ|���?��J#�H.��Q��O� ��n���l�2�(�4���r ?���lbm4��3:�N��o���*���ȋi- xu�}Lo"%��~�Vqe��K����0*�j�y��2�ǉ6� ��a(�_�J.ݔ���W*����kB-Ʒj'�i\�{_ש�<�J8
�ɞ���Rs
H���8�SRo�WWL����4y�������a��e�u���S�}/wPu�[`�x���$쒅t�L3�
�?��o�b�.8 v�nm1��?��,[�i���i��]�/G���9g�<�stQ>(h�<�qh��4�����e�Q�>
*��u���'t�2Ȧ�h��\E:hS"��_@�����~���F`=C1�o7�S�h85:qdUC�u�h؛�� >�����x���n�s��b��>(h!�kQ��۵	|��:-�
�ʝ�z������%��#�+�CG4
�^�ж�>�q<����}Z\*��m��ڦ J�Jv������)	����Ѐ���Ʒ�$�o8��øa��1��V_��рL��m����1�g��L��"b��n�F ��F��� ݜ�`g1�[Yu�;�����ˇ�2L$�j5�ۈ�>�-��(�����V�K���U����^K�3.���ht�v2�����毇��c|�� ���j�� AOS����"I�QF�h���B;&�>51�dz�,1� �P�@��R2�L�ޞ������߈�d�^���Q�!E�o�ґ��c���ճƯ���Y�v��8�i�х�1���fM�K}6�.ze�ef+"<�E����u]�U�qșŉ��ȳ_H�Pg� �b�W0�ű�DR�4�X��$GN�Б߱�+�L�q|��V�p=�C�s�8�������㤍��O�KLef��0_��JySd F�s?|��_@$8q��J+�&G��5�ǽ�~��rK%uSR�U�1w��5�=���~�#͆H8>�������(��[��3(S�n^8�>m�����-��%���4���Kf�k��t�ЕW+6c����C�-��*�"Bz�>��z�O�0��c�%�s��2��ʺ���#�z��VK�L�×Ź�x�XS���+X�>d�M����/��W��Ư��:�q�xӗI�`�䲧�R���"b�2le_��`��NK�6X�C�.{^��3��ݎKWs�	�ÚR�FV��@��{H�͉��w9��I̊�ۧ[g2��S��ɲ ��l���6�0Z���Z�ۓ�'Bvh��١��J��SV~K���t����B�J�,��}��&鵲�B>�څ���Ϝ�,�pO��f�m��?��n*�""X�WAU�`�J�N��_K�p��7����/>��>乪X�B´�a���<�;���tT�!'r�(��"���(~Y*�l��W��Q^�p�?X���|@��?4eg�1�=1����Ӝ�g�*���g�l�yP�HNx m4E�B�f�M���s[]Ж�9Q�1�Ql��@���Uk���2~S���ḷ�:uF|���:La���D�!D�J�g�#؜���NT����e(O���	33��
�.A�^�nN�L*��Bm�|���j%���E�E�
B��x�MH�вI�@�"̝��K�&��Q�	Ig��u\��H���?���g$D��W{�L\	g�1YD�%n�9�ٰ
� K��2ҭҥxȌ����d���2s��׋sÏ������q�`�)�m{T3�z���/_J��K�1-8!�i��F-Q�;:L���8\��P˨}�ɜf�QAFn?���[�۠\�F�~��/���Ñ�O�nC���� v�C�ք�d��'H�����ILυe�]/ȡ��k�[SZ���:#�Rd1��TU���¬��WZLb�Oo��!n�H�߾(+�M�GCS���r�T �e��B�/P���y�_���3���T�W�?PZH����jV�Ҵ����K� @�z��v���'�Ptj�&{�X�Ԧ�.�K��?��L�)NM�������b�@���3��*�d�s@肤v�A����b7�eb��UD~�-�,,D'��6^��2�s�Ҽ�������X������	� r�x���E�;)�k1yg/�PUWSF��Ԯ�od!~�;aZ_�h>r�� x�qc�E��E�ʂ�붘��	�*�pE�K�[Z�t;�1���aѻD8�eC\���>/-���d _�Ŭ�OѠ���w�v�~e4��i"�{��~Wj/�!����LI"=���h<�17��2aU2U8� �R�+�����.����4b0��F9@��_�N�:��@�g>m�s+��Z�#�g#e[��{���9���}'��Lm�¿2� �U籪R5�ll��sx�He���/d�����%�_�o%����0���ⵢL�����4����=B���{2-x8 ?��u�/�/Q`W��a7�U��f�˟����Ok�dqf)_��A޿���$s�}1%�K�_�����NMB=�R��'��4w&e���i���6��|�JV@hj���D���!��`ޏ�K�z�[�zoMHZ/ L�g�ʲ+� �&�/1��;��aBkˍ7�rA���!/J^��E�z��j�g�9ͭ��Hm{�㳰1y��^�E��Hl����rr�f9��Xh��ܣ8�d�;_����D��Q������k�aNV� �rк�N��OD�H��p��+�HO���L�X���1��ٸq5Yi{�zp<�:;��A]��c,��@~a�j@��d�/�Ή(l����fQ��~���z��s���7�N�	��5\2����;�k-Z�Pڨ�d��7q\Cު�1�eur�a4���W�p����NFg���\(W��]C��#��p-���g��#��o�|�c1|�K�OO �������B�]%�&ګ���*ye�4?�3}�%�8�l��ڶ����#6���&�Q�s ��OL�7ȏ[�i	�~����=���و�h�� �YX�j�[���w��2������K��N�B�v��*����~�o_�n�*Qm�Ǚ��!��ht���[L�T�]M�e�~��繍����LsG$�3K������ﺌ&�EOEd�;����ˎY��l�]MlO��$sX�F��G��"�(7���.���+q;��@��6Y��P��Њ����*�ہy1˜3���-kaG�\k�Vj�p�ɡR�F+���C�7m�_��B��ۊY@4Gh!��GV˃�k
�&v�^Л;�-9�B�~ӣ�X�dө���P�4�aƤ����B��"��rU�H��e�sE�a{j�X�ş�%R؊)`�l]q���t8.ٽ�Wm�l~���e��H&3�m�l���#�h0�_���D�)�[�9�˷᭟$��Q �i�(��5��w�/)���#Z�yW�˞g�=���]��h��2�C�q���<�����
uܸ˿�f�rSM��vP�<���qq������x�x�O�%��2�3�{q(�1�e~�����v���d*����B�N��|6�I�s�3�L2&J�{��%�}������)������[�\��lUu8�z��8�+��h�:=|��s��\-ï#<ʊ�Ղo��F:���i�5B�K�,��jj�=�^Wz�4^��<xgsQi󮯈�D�����6 ��@$� 
q�N��&	��f�e�q>]S�ɑA���ȵp-��j�D0�6�c]>'Y
�g)��;V>���~�ǅ;HhҊ����NL\xH&UXA[�a�#��:
ę˻;=�؟�xrK8v�P�X��ȞA�����z{Va��g�N�2��Y{A�`���4�b�s`�����/��v�Z�;�ϙzie��	�lz)j�q�.Ek�q��O��V�Bn�o��ΝZ�	H�l]T��b����������1����6w��&�$�'�'!�
3���呖e�ZPT���n������a��?9��z��`���NUpJ�jF��w0���U�!�K�����J� <��ڂ���ս^���h�+���P���pZ�|v��V�Q�D�*"�ф�u�J�sS��985���֞��=i���.?g�%�E9� ��I�^2���!�|����g��eV�$�Y�Y��%%ȚS�v��О-Wן�kWR{���E=N�%.Ìǐ]��_<���a�ab�#>i�v�[1��9�gC�0JvQ���-����s����,c�\����t�D�����'��@L;V�h����p�ؚp��"f��t<�[��-xI��L���'m�^��a{ld	l�L~�o�+n�=<s+2�+N <�zFe�p���L���ᣴ��3�����F���W%9}r|� >�葿�֤qa�i4d��$�r�ǕMz�U��H�g�.��!e�����M�:e��U�{���|��6�i���{�ܣα~�J�\�%���]��^{jBBc�o�`�z�{wN��r%�k&�P8a���KL��|��'��	���y�J���~��V����B����ؗU.U�35$����`�]ӪHdv� 5�E#�P- o���A"sR��K���l�ej��lk	LN;i)��g<.��YE��$�I�/
�ҥȨ.b�0a�Z�6z�E�k_?��߷'9��d����p��"_�B�"��%������������)��T�Q��������-&��H|p�cq�,�r�#�O�x��\����eA�r�����i�{/��,��0"��$�v�;P%�Mp~K�>�L��2���#�Ce|�e�!�:�Ŗ�ERg!����"U������ҧP���O�:��Z��2cgB
�=\{��[	�b$Cp���׼Z��\��w��|22�@߱��Џݮ��N���	Ծ��ٛ�����5�z=�����}q)��,�%Y��s�@RiG��{MEv^ }������&�A���b|�K�\�pȍ�kP���O�y������FbJ5��E(�c�z���Zx[}���%���4x�ZϘXb�.��IuQJ:o�qȹ�H��q%�>��pWGF�#5i�w���"������|��]-���7���
p�m?�zDƨ@�m�VЃbΘJ�Lq�P�:B���^�/R�XL��3QB!�ًL����|R�zQ�<6Ӈ2�#`	Q�P�ّ���r1b��9���������V��F�=��-��F��H�z�������Q�@��I�~���U�`U*��Ro >T��D\���<"M�Wq�sy��M�	��j�}����`XATy�<=ō5DZ��tZ��|�Pk�=�Kp�lS6Kg�M��q�`q�m$[cP��u��e0�k�E�6�b8�	��au��"�8\	滄�x��.5�h��)�D�t��R��#1ԟ�D�b�� ����B�?��2��20{7�C3F��C5�I0� 澯���� ��L'Q��V
�g� �m�b��%7Q0�(�6S,���5y��%ÎI���F�~��X����*iH.B3-�X�wj��woc(n �g�J�eR�;�;�6�!�沼�҅�t�+ <
Uj��ne+�~��R��cz���I"��byer�>zW{]D�Aش�G�d;e%�o��)�Y��:�1ER�-#�[>_����d�	ЯՓ9ݟ��N.G�W ���zv���D�	X+�s����V���C�і���	+2� ��4���V���m��U^�JXom�N焺���p�J+�����!}��g��@�)*װ&Sh�[�S
ׇ�h�S�$�U��E��x�*�mJ�&��OZ��`��z�e]�۟�nj�h�.�ݾ���|���:^\Xh��i�.|�l�OÐ7��{����r��ۛ��7�j�Q�Ø5����?*���D��(ҟP�-��K9atT�(#!oj�s}$5Df�Rs}���^�E�4<�"�~s�SK����2���������	��/�>l�j�x��7��6[��,��N�N:�q;V�/��1A?��Tv��HEFAǀC�wQ�@���[��]���v��jr|�4��N>&��\(��2�(���?���GmN�V5��\\��;�x
<d�O�����	�U2�n��OR��z+�~���08�� K����u�e����Hi��ܱ�m�P�ZܳUɉ��/�{��@����
0�mWd�(P�ɱ���9l"��S�#���Sl7תX5؄��"软�تD�Ԡhď���Pmغl�5 ���V�����@`m�$�S>x�kj���K����W��n�Z�T":ln�!���E�s��v9�P��0��誒�nd��H-�o��n�1<D�"��#x�:G]��b��L�6�;)3�~�6������J�@�̟t��ڷ��o�n['�%��Áb�,��9������w�TY�b��	����yTFKSZ���F��hr�2L��T��- rD�T���Y���<��ﴠ������1��~I"{�8x���k�����j{�BΞvW��� ,(�<�э6���؁p2��(6q��L��["�u����C94��
]�3a�]1-Dr�Gě
T�~+��ܣ����,5���"3�-��i�q=���p�DX�Np��?��5(!���4N\΅�ߙ�4�v
q���!�ǳ����6<��<=�jO�H�`+����P��Nэ�j���;�G��CT�}�s�
H�Y�Z2�4. �߽�P��A�QP�k�c	w�ɻ=��.���n���!����!����[L�3;�.-�`�}��;�]sQh����A�S��v�j�>�}�Α1^B�d����H�q8R,:�������_�r%=�lK���WڵL�e��{��C���2��)�7��]b��E�V~ۆ�F��H1��ϡ}(�$<��7|&��[��Ԑ�:��~<i�4;]�&lE��~�7:hN��'��rZ�> Ǝa��if)����<+������D��*�B%���=�V,i��������a��T�r����,A�4��c����ȋ:3�i*��6�v�E��Pz���Uf�%ˋz��a\���n��/�PD�)K=�p �cƈ�e��0�RvQ�~D= ��P>��܁'O)W��*�@Qs
���}� ]�ܙZ*j:ef]L�Z��GK-}���7}�u (�z83�+0��4'��{W�o^�!>Gb�b�z7\�ָB5s��J��۫n�ݞ6�X|����^jXԝ���ӹ��2�\)_�GQ?�Q��ap�sR�C�=k�d�i�e��V�P��kZ�� /��QL`��U'hJ[i,&6�owA���ߎ�p�[�'��������!
ħ�0L���Ԟo<�+��㛭0�a����w�����[�m��Z�	�o#b,<Jޛ_R�	�ŞE/��m������`��c�<{�X�X��fAQ�p�ʵQ️��Ԍ)]�X~6�i��_��qS�ڕ�1%�P]��P�bŞJ�חf���@�yG��v��(���Id��V9�W� `�9��c8���Z�T��>j-���(�Z8��~�q��ő$�c���l������۱���N,E�&�����$�8��j( �� >Oa4�� ��>�ߝ���{�sT�'���%󺺧��" �`�zF=�^�S��䠲`�����W�Pj�������@�sZo$mD��iI\�iA����7�SW��#nS�Xɜ��'6�X-IU)��[��tf���)�d̽2�Hl�
�!���żYQS���p9�-C;+���pu��6�]3W�*�8�k��`̱dŗ�,��Z��BF]�{0i�#�sb(}�@^qW] P���ߋ�dѓ�	��G��{v���|&�uK�nڔ��W�+�/�پL��;%q}��$:`�I�󼟔Q�����c��WJ9<�8�d$��}i�r��_^ߣ�y�������zO@Jj4�<Z�뛢��Z�=|
X&4��_�(��@!,��9sn�/e���ғ�;���F^^�bqDϟL�E�|?!���4rU��f��3W>�Zg^{w�G�����x.��0(�yY��!vJ��d)(߼z#7v���]���hsXM��_��<��mO���������#�u�Z0��Y���h?����|#1x��@�8�����bނb�Z�&U�A֩��Bs���j���y���C�	������Ӟ�Yȓ��<x��[�1W|��}��B���G�AbX�sϟH���i�
B� >�SC�_�,�w�w�3�)D���JeL�}�o�bH���b�miG��Y�To([9P�t�6r�=?�ORo�Jo!HK�P�!�Q����SNo�����B�*�v��1u�s���r��E���jݪ�8D��xv"���]M���P�sA�%Ey�&ࠬa�<a5�7��ig#9s�o0��}j/{=V0��/���Հc��ey���7ăO?�Nri��t5H~0/�f�U�������_I��-�҅�\u�p�J����I�f+?�����>�r9L��?���n���~�S����D)�ah��#���YZd���.�e�ƹ�@M$�A��Я\)-Ro�i6��L���B���6@c���o$T��&ٵ
x��GpF�k�/�^���	����N����ٴ��L�Ҁ�prkK��HD"G�vI���O���q�eMJ<X`������]�©�}�����V{8�<���7�pv$��0����%)$�z�4X�xG�㠢�� 
�����3�d�>�ud��hG���
�l]`��:�)�4��]GFgȺ�xE`.>T� \�ǋ㱤��P	�Gg�G����$r�1�2�<ֹN���i%�?�2��:��7E��H3��B U-}���+a�#���W��X�{C�����o�7�=�]�rP��D�J��!�\�h��vm�?�ԃ���ڰ��ۚ�5�H�'�M�5���V��ݪ�Ĕ��}X���*��;=7���WX}�'O��X��L`?~�c��g�����1csw��D�1xa�F�n,��e����!�1����M����8��E�����x��J�s{��!o�U����2���a�m�]�̞��:�l�m�@���f�KZ�	qOjf=DG������S��A
��s�������?�G��qT��b\�Z���P~�����ß�-��SLɫ�8X��1�鏹R��f�rܩ�7.A��[�' �#y�fm��@�yf7�su�ӡ�g��K�/YϞ���d��f��}ڼ���c�B��I�$޶��;��v.��Y8;(RI� ���Woz�0�)��=lJ���lu "4\�%�������r�����&�;�`4��nzc�^&�����f��m����K�M8�=��9�Z��c$��G��Ը91���Q�k o�y�yR$<��S��~�b%D����Cc����o�J�}3=��6kI%��P������d�{_��5��14?%֑�0�z�de��6��A��msE����\�ё`�m���2JR�p�e7
��'�!��f�&;#\����$B���n���ׂ��[�������H����W��Ǡ����LI�CC��p��,g��[`_�#8����i�OT���������F���0F�0\3�Y���o��>U)�cgG:/�m�^6w�S�]�x��3����:GЬ�N�!�T�����ը�b��"i���p�,�7BP�kꏵ�+��
_�A!WA�3xzӁok܉�7��0e�R!�`[[U�&���Vq�Y9�D���s��_�r�rD�R~>��62"�:��_ָj�����F�Lֺ���|����'؈�v*J�ӓXG����G�o��D{�F��W�d�!���n?ǉMX��H��Nl�����@����wS%�D�ɝ�@�����"��A��ܓ�So�=��|�j�p���YX����Y��AyC��&��Oō�=�)����$���I�ࠧ\�5��~C��`m�I��έ½� �n�A���k�'4+��^ ���A�~��Z0�*�V��z��rq�D�{�
ɖ���ѭs�n	���tE�G�ē�:��Qi/���W���㭟��<Is[[�Uzl�b��:�"sv���O�KwA{����^�(&����B»��B�͟K7l������:�n`�M�>S7O��Y_0Ϊ<r�� %���A��$b��=���]��g'�ʓ�C�JF��EPK�NQlFo/N�a�����$��n��ѓf�=�l,:���F�^6����peor҅�s8P9��^,�Xeڕ	������&����A��n�Y�����3�!p�h�i�XD����f>/�k� ��_C�uKn���(�@H¿���E�'�Ե���3O�ޭ��`��A�@Q�zo��-:�����9�P9����
�@�!� ����jGZ�*%Y"o�z'�Xp'�Xn��K���a�~����n���=.ִk���pt���E���N%�/��2�u�(��/tj)g��v{��s)�_[@T/X��h8L��@�	��ԎK�N���D5K1�ỳM�뙏�^��=2�j�Sz�jw�p���Q��� N��.�ć,1m9�"�!2E�D��W���]��R�(JR���(	(��R�挿pB�B�'�Sv���Q;���T#�Λ��zw�ǱC`�M6*��J�B���Nk ��`����T��`0��F&���]:�+����:���&H���y�$���V\Z���L��1__�����0L���u��C��K�A2��UL�ɫ�flR/g)�3D�善�q�f�VdWռ��U���x�?y���(^�GwY0;���CF��glJ9-,(h<�i1&�[�K:m�B9&��q��z��X��=���'�T�"��9���RB�ΔG�Gt�J��;��܇!qNajR4�$'3�����O��{^�욎 p��/�(�2�Ѓ�=��>����  4��{Jϖuk��w� Ğ�0FX�;	X�����S�D�����qZ��C��e�8P�}4��^>BJڢm���'�0�CI�z�8��-��m�&o��Ұ��͢��:��~�����D���������냋�a�"��*���W&��Z�@�����I`"�/^��Uzи�ߘ�����__0e�|*����\;��<�ff`k�U�	�J�f�YF����D5L^�^6#$��t��
�B2��E��~ �:���������5���P3��a�Sz2tƜݏ܆A2��$�	��~�?�9�W b��w�IL�\
���D����L�Tj�e�PV	�ms���!8��WR|G�?���A�\���/EG@��JKK10'�t�`������%�N׸e��((9	=p�q�c_7Ҟ�Ynj���Wrm����-���"�F�ђNK<Ij���Di���c�^�Z��?�����+m�ҍrm�K���Wh��Z��-�=�F��2�l��T����S�!�R������b,}�*�0���f�俺���p�M���c%2�o�mϐ�ܽ �ZW�܅��v��eγ��֣�E8��
�b��5��Ѱ�Y#ܙ"��8��R�)۬0��N�ڜ�B��1/����2Rq��Mv�o�+{/e �&˲2��*_�����D������S鮫�/�jL�Cl|��vi�1���3s�@���37wm���"�C������?�����+�
[�x��U��Zk�Q�,.��iK�|�s9��S��@��Ag�?�8$E�]Jv����)#AЊH��L�̬ϲg�� 7򦩒Ưꐩ�O�ҍm�Ê8
�
r���n�R�5d��!&�YF�	 ��48�S���'%�=IE�����ɆƯʠg��já��p��6�Eю7��c�'\�oU��+p���g`SM���y�e(� �Y���;M�cp覲��Y�z��5�^6X2'����+��3]�m˕7㽪��G����N�IUR��J����`��t=ߟդ��V�N����8~�|��-x_��=�Ҫ��'8.�J����w�WB���!i����ca�L2�b��"�+����i,f>�y�ً��bF�d^!L��a`�yi��f���i4��O�Iŝ���<Up@����	:���/r�2��#߫��U<�&���A$4��*�#�R8��q�q�r�Y���|�CƢ����i��(�d�/�.BW��S-o��ԯ��?�� �w����ƙ�t��<�aB�`�Ҵ-�G�&�%$��{�'��.��\J��]IX�Z-CE������`�}�3/!�ڗLvB��>�N�!+�?���lfx}����PK��cX A%2���e<?�h��.�_�A��%�4߯��*�Z!Ѕ��Xq?7��+^HD�����TY7����]��BLi!S����B�;E���_�8"�?��Y�K0����yF���s^?�Hc@Z�y����+&���+�_V_�Y=&$�LO䂂�\��)v�{V-/��&�v�h?���9Փ�/g�a�j�c�l�;�$W6X�2���|��J�v2�c�MJE�n�,�Cy�׿9Z�J��I���AP�?M���5�_V?�{�τ�'���@Y!*{kj��9����- �_��C���Q>[��@o��@߭�z�O�#c���	��ɴϦbHF#�)�a�kN�Nv��n�ٜ8q��J$hF!pW�ש��[��	PKK��b���bG�b�i=�gt���4��A,�Lzy9�-ʓ��Bsk���^���U�!.Њ\�r��7�I *�i��� n��8v�R�hhVU�ۇe�+}hU��/� �@4�"1�%�%]M�H�b7U�mq{|�6ۆ�ii��(	<Y�Ť�c�\��.#���T>�^�$�6ԡ�*�NWg��Y��P���& �zN���O�*Ln�y�/2C�Cc��p�	|U�>\
�G+�^g�����jp���U����u9�YJ��s�Eizm�r-�̽x��9�Ş�+�V�J��9)�m)L�ON4��/�Ci��l*�A�oS��x�5jf��K��}�@�|����U'%5�9�J�W|\�H�`H�b�^�|�� z�_#�'�gZ���5�½}�Rx,�b�����yw���rGr@l�p��l� ���w��i*t9B\F�U�:>�L�G��I�JX�M`f~2��`�d'Wa7��p���\���|�gq��C_���8�X���I[tǝ��ag�8[�Ɠ����U	q���Y�VCm Iqh���x5���B���X�b�^�Ub����!�w:1�M:ڝ�&ǥou�by�~,�# ��X�{�Y缀 ��_�ҋ����l��ٷ}�oz��lb���
�Xv{1"�Ĵ|�S(��do�B�>�@$0>�K�Kla�^k�I�(��)һ�g�WF�|
����[�&�$�ǂ#� r��y��T*
d�
�[i��1�`5aE��|�T+�Q�f4���B�����M��l~K�:IWdy&>D=6i��|/5T x"%��6h�/q3��ٝ��B�,�vۚ1W��}�,c��Z����#fS*�!�-(�P|�!�3�#)�O�U٦�����a���d��=U�Ӄ���;�h�N#����A4�{e7˭O���.-p,�yZ���)y=tw��/��ᡸ��߅�*�IC��ڛA����1���@��Wg�P1֞�������Lf�����+���q�1��j��/�;w{�Իgc�����O��m�}`Gy��ٿ{�t|�Is��O��cg����F'�i����^���~C��.pw=�!�6y��:�D�u)3=W&0��|�gk,|��r�U��3ٟ���+�n�о�q�?�����[�ᓂ'�/���)���?���C\����6T{X���z�	����÷��������p?$N7�<���lS�K;��� �}�������)�����Ӹ6��;�4����١�o����xT��xGH&���ᜂ�3O2s�Sc�}��}pu'��	*�{V��7*(�J7W���'Z6�@�+P��~{�s�/yt:�Z^���
G/�3,����0��؞��z�e���P��v�.d�뺄-Yr_��!��>��o8�9����=f�q��1����>������2�\��2ě��.�~H�|�y�spl�fl�S�$5�����K�.Hp^p�3�P���@���8|q�:��#ff��#�������9ikWy��X�^��E?m��u=J]ק0Z�}�U�ur�r:Z��-_%!G$Q��ߤ!u�MX�$�`�9�Q���:h,����J�}K�E��D8�LP k,0���4ˎ���J���?�A!�{�w�.�=��6�b�DM��P8Y�0'�מH�:�t���bX�Y�ۑ���/�+��gǟ@���Ϸ�h2�E��֛o4�b(�����c�+^���(�M�"���k����@���A�T,�.��-O�F
��}kO�|�K���:Uh���|O�\�8^V< �8���]n����CxUP��st��7�í�)�?��ƧI��'������!�C�w"�v���6��,'`U���Φ�V_l\N�?A䪕�rx��ǅ��$����H�fS �����Nc�4$�Zآ> ���qR��ܜ��@m7�'a(�Ɠ+��$�er]tu
�G���9	�ԗߑb�����t���;��Q�쟛�R~�(�c���!l���ޭ;<�K���mZYC�W���#$J&��;y�Up����$���i�T�{V_��,Sۦ���!��c�m3N��� @<�?-��$�}������G�]�JNע̬ !;*F`��h0�c�7����U?~��a���؅�1���q�dBv��S���S-��R r�dy�����Wޏ���V�xtØ^�*����^�^���J�l`Ig^��<!v�>�	���^uv����k�C��o����]���	���}���n�7޻�cV�!���ƪY�[��|2�U"�,���F�A�?a"'aRo�C'�����/�k���# ��8f����0�=���8;}��Hu�ђ�N\	�/8����Ʋ�c�aj"&c;x�஬o�We���;8��g����qG�~RJP�T�p�����m���+��Y���������ǯϏ%����+Y���f��Qj�:n)�|����b�@��jy��_h*2���������]&��H��F��/�m`Z�F��*0�2�[�~x)WU�I�?�X$3���^��T�yK!�7A��B�Pϒ���Bg�؂�*Y�+�DՖ�� ��ٌ�0�"�PJIS�<����@:��`6h�u���G�Ĝ
��|.܅;Fq�|�gN�;g��f�oC��}�Ɩ]� >B���< ��}To��n�޲7e/�����xۦV\�D��>9�@v���%��{���y��O:��
�U"f�szC/#�;�$u�<nr��
$�eq���xm�[�f:O��)fY��AۀԐ��|x��>$&��O����f��	@�!�)��>��0*}Ob�z��@(Ϲ.8(ۅ�{�jf;�I�H<�f���6(*�}	C��P5y�(�*;�͐�Bd�<�^šՃ���O�VG6Oᕆ<35�9oZ,�"��7��G&��A#�bY���-ts_(��.?{�pd1��ñV���>�¥)�m��y��i��7����h���V ��g�v�_F=�CҜ�a�pV��	cc��5C� B�k���4z����_���]n�>}���ӌ<Q��ؕ�J��y�֘�~�F��sI9�c���&^M��_���h,P�8��&�H���Tm�kD�-�5.\����?uRM'A	,�l�1uNC�x�c�>��E9���8���?��6�5"��z���A:>�N���*I~����Q�Y� Q7�ڸ�s�F��._N@?h	w�T����%[��U%9�
��^�P�F/�a�7Pz��L��9D``n���θ�����)VS5��󟱮�WW�yc�J��W�6�|�,��"����a���<Mf��������0���ň0��.p>{���V2+ �wr�ei����M^c��j�����e��2��ұ�T]T�P�e?�ʫyjN�@�9��ۜj-�p��A;����e��j/��4^��w��!��`T��#��� J��z���^� �i?�T�I��#�K��XH]�U������ѣ��&���`x\�������y�xUuVTj3ё�F:�l��Vw�F�=z�fqr�k������Gp5�m�/�WY���vr=����9BG	�m�sz��$���5bl�G9���b�{%���)0�:�I�����<���t1�������@�����ЈZ�����4��#��� K��]�{������p��a^����*q)\�y?����;��o�7�FǇ��҃��d�P�e���|z'W�&��?,c�Lkf��0�/@bE��k*�y �a`XL$0�	?���/=���ҹP9I�����m�����j 16��&�Q~K���_y����lf���@J3�3�N���D8��E��ȁik�R��0\�?]!��;���/�N��0�CN���T�j��J5O�`�t��9��֫w��/�&H�������`�Ht�����O�N��	�"U�2"�?�P��݄ܻ�I���� m�^�͂�r�]1{`�E�y�.���ĸ�Z����r�c�;w�ä�^�5��r��:��}��I��?�rtڬ��JT���y ��<�k��ckZ!t��ɥϯ�w����Ti5}]Ǐ9��
�p[���U%�e$A#=&-Vw�|�sӺ�潗3�^����x�K�XaU&����C{@�B��0��G�p�iB������y�]*?asz���E"m]\�߸���$�����5�����Q�<v��d��ﶜ�|��x�hl,�7`Ї	��"-T���Y���
S>��PDm3hq֙��a���@V�	Р��}eƇ���;���fma�8V��HM��Mx�@�q�.&��JIyP�ι���R���3�ч`R��W�6'z7q�M��ac��&��#�}�I����hv��v����;���m�M�D��>��`dC!�aH��.s�E��~u�ַp͂"(M��}�!MPW�{j�Fxn_�I'M�'a�4<���l%�=Љ���rO��*G���i���z_N��/�����Gkˆ,��R�ב z����t��7y5��	�jώ·�^�'�q6`�,T�V��8q�U<�oщ�&�"h���՚g[=������TN�~SI��U�,[�|�H�v��3
�����1מh�����:���'P�F\H˙�o|�p|!y���ѣ*�����`�aV���$=w�P~R���7�(�wn`�	��ڶ�Zk��Q�[fz�eY��Tx�ј�l���@��9̜Xhu!t7g����I��M�x��e�6���l�fy��N ����.�^�٘^Tz7������\�tʏ=V	���{�[������mr�T�"� ��6��47���f��'�F؏V�scHN����Ngs����D��Ș��}��Q��="���s�Ȕ><����ѷ%/<~�����1m�;�e�g�2>�Ir&Z������#|"�f��?N��K������?�[P�GI�o�#� =S<򌓦 m� d,x5��l2�eI�j�濣��ʄ��N�q�D+JR��{'S�x�J�u��5=-��C�~H�L���>uu�$��5��dj���o@�^;I(����ǭ����xo��Qͣ�p�Ts�[n2�x��M���wH%�2K&�V���?��=C��U	\Hzv��'�1��iH�߫��mG�?�	�l�����M��?@b���
z>*1z�˼d+��qWo��ϑ�cg(�9��e�^X�B}�,5�E�rJ��R��`��vT��qY�}ܥ�
�xLA�Ϣ��Ѭ���[P7���TV��c������1�n�W�w��i�v��?0Z��R�x�׼U�R�w�8l��@���EP+����^y`0e=�#JB�c'7�X����J~p�I�[1O�m7�O1Ju�c���-K/W�Y� �Ѵ ���:�U��]`��Y�����%�VUy(^��b,�9��(��&�3�\C��ZM�D}�&No�0*�wZ-�|(
X�C���{���۲$ڡ:`��Fkæf��������4D8Vo���o ��6z�.SS��º�)3�د<�Kf������3�ƨ��,��~���7���x�6���z��c���n�! �h�4�����Տ8Q�+>6���حi���,QA��%�F���٪��x���]A�H8hĿ��{���Ĥ�ym��J�^ݪxk{����;�\ ��W46n'&��Z���s���tBl�0�xq��q[��+:��s@��dUg���� �C��ܳ�C����^0:��~��r�^����16��@A����Ajl��Ղ��k����p��=kD�M��d ʻ�KM���a�������B�YvZ�r;�\Sy��卶�L>��;[��Ι�djh�[��T�pB�e����&�{�������~K�8���j9+CN�;�������[�
�{ �d\�v��E�=Ry������Z
�-?r�r{�c�3�c��j��,��b;�E�r�)[��n�},ǩ�,�K�ׄ�E�}Ŕ�g��&ز(��;���1�t�
��K��/ͷg�b�۵w?{4�">�����Iu�*xǋ ������َ�v �L���}�����1�c�AgS�97�7�hg��T��&{"t�:��<�;�M �߭��?���K�' *�L:q��c��M�ݓ�X(k�}HGީ��4���4�ڪ�(`���6,{�ΫѰ�TT��D�&5���g�\�sh����U���Spr^��O\ښ�d����L�t;]�V����f���%z����Oh㮭���ʃ$��]%�̸kbK�y�-�,��\�{v�@�?��ߡ��iV�4w�B��g
���lo�-i�>�S64͹�=Y�М�4KQ
���{���)�b��O���Ӗ��)�%]���v{�\1]LR&��������u���	�C[�X�gK��¾�%��� �闑�����%��D��K��X�.�����d���E�O!�)�2s����H_
��S*om(	���%'�����.��(�S����������ex/IH�����O�@�����WB��(��r�*�y0��Z����&ܸ��ֈi�z$��&���>�܏�GK$��r3�{�6K�T&O�_i�7]P�>p(�}Ri1� P���u�*@Ď��d��Byh L
���	��"��ڦV������2���P�Y0*�s��N*�E<v����t���"*t%]�FԮ���Rn��3	9uz�+���Se��u�Co��;	�+e������*�8��X\>��=�iI�΋j[QR1�%U��aQ���g�I�K٧ D�s��U��9�z?"y�z�͍�md����]�9Q� �=��\��V��i���#��~���&V�~UYr3sx�~gO��N`��lٗ&+�C��h�����ϰM{��)��,QB_p���.0=k~c�$�NE�}a��r�^��?r�<��1��3�i!s�U�����i�$��t	�O�6ٓ�}^%���^(QBS� :1�۽�Ap�����dup���d��T�VM�e%��T����V7ɵ'�������k�uj�e}���#��!]�3�;����88��u��5){�)?dxu��b���a]i����������̚�>]O��[��a�ݍ�|�c��[#+��Jߺ�� �y.��|劃���fM��ג��,}�T{�%�5�F�o`#3�{�O3iZ}���nt�����n�E�\���VR���\~��� �P��3&��v����N[z��q$�J���i/D3q�-0���{{�G�bh�d���G07����(TR�υ6*'��l��ے�?��L��J���[�uĥ�&��K���C����D��؏r��䬯e��8�_K� �=`�� �����S41��%�0��nK��B1���V��-^�ߩ���#&�����m�TD��0���n�tE3J�y`y��]���e���m���	�R��X�Q4����G����% l�����}[�h�)PX&O�X�+�<C��y�@������v��B;��]��Ճ��X���d�(5
��2r �����`(X���L�w���ɤ�E� '�w�;B�J̀��V��"J�8�D�I:c�# �2Yn����v��)��Dl+p��Dӽ)�6
�gJ-踇ޜ9w�Ko�D<�C��Q\e#�Ѧ�	��n8ɯ���>�N�(��Ć��_�}^�LfF(G�S��;,�����.ը[�f�KW �(�S�h�OٲA7��-�\�^�v�xV�?ή��Mפ���A��5e�a��}Ą���Q0�QGR_O��tc39VQ�,+�#�r�Ke\h{�2�'"y}zR%[+�y��[����Sw~��{.��p
f�q�~O��?�����(ڟ�x�'�Y�C��I����J�b�g�u!���zH�(�ئ�?S��XꝊ�W'S��C�r"�X��9��G�)+?�X:��6}%�de�i�b|-@Wu��.��D2�>R�v|P^]�f�I�-���Q�m �?���b^iocG��NoRx���:�ׂ���$z�`��݆f��=-��� �m5$�r�bR饡<	):9���K@�Hs����B��XIK~���H�2�e.�4�����Kbo��6�h*J#�[��VO4�,QJ��u�r����i��$0o�^��h�@��k���o�jۿDU�X8Oq@�
�4���ߊ�����*�͓����R0��6
�4��X�r]U��z��e}\�+\?�!���6�N346���1� L"X��EUW]��y��O㢨���>
 �W��4�>�#�֟��"�1�� �Vb���7�.��T`3��ېX��9N���<W<�SS��vQq0�_��Svf�1����"���C]��n�ؙY��v	C�X�������Ye�������S��\6��Y�������?�K�ִ����OS��Z��~�
�k.v:\R��A�u>}�/�d�KdSVu!�4��,�u�w6v�"��W?8}��y���(���%�ļ��G��܉.1�3��Tr�G����������K�hx.rw��i�B	%L/�n�n"��f��ݤ��R�E�2��:���	�7<�=��x�����u��-�a�����D%Q�=��aw�9�M��@

�����^��`����4���c��!Ν�|9
������w^�?�ƶ��5�l����/���@���A߃/�ݮС4Z��S�©	oHZ h �Ҫ��yZ�Wצ�V`Z� Y8��c�E����c������_�HSs���|>F���o����+�ӫO��V�S�I�Tkj�n��>);��}��n���}�A�T~u!t�x���9�j���~����	K'nHp:�U	{����(n..fQ���_KVE�}�3�&�˯Ho��>�K�R��v��͖��\��_�܇=;�	�E���^�o��Q4�z�� �"��gW	Bh��K+ٯ@���� �< ���w��Tj �k%���+��~g!ĭ�_��F�c�9���=$�#<�69|H�ѱ�����뿅�'=�L6�I�l�c6����.�y���Y��Y̎g���+h�*u�̳�X"�X�,�[)X:4���5q=asx���"BN���mz�0Ci�<�^q��G:����?xz�"�N�S*{��O.�.
 ?\�6A�KR��
e��u� `v\mUJn4��a�4���?���r8Q�k�����[0s��I�U��
���<֙EEq�>	h��N��D�@�#okN6�-x�˝�L{���Cv��}�C�C���S����f�2�H���e�+��k.�sM"��[/��"K��m�@KF������m�E�^4 �\��d�;�+��N��Q��|��v��y!��B���)L0W_~l�ք9"g�G���͓0=�vQiZi|��	��q�1���Bh�B� ��X�x�|]H�FB�D�� �Z��`��L�֬���i�H	Y�>h#�W)��(�%�n�4�~�hC�r8�Y���,�=�T���mNHQQ���P# �u �v�E�=�VJ�@��gv1i�8
�n�oD�e��d��i��.M��Θ�H�"=HY�6g��Q����u����4 ��j4^�ʄ�VvqN�����	/Ӫ�aH}*sY��ؗz��'�b��r�|=���;ͣu�r�T��6�������U?�C���Ӻ]�q�#]Xg�uY%\3h��+���8'��Q�q��g&Cߔ�����[���5��)j�H�0Qz�FFq��q��}�UH"�`����j١E������Gs�Ӗ�׉�n�u�@i��� �m�Y�1�S�uob�Vh�跒��F�N�E��͕+kD�Ї��o�Z%ut���h�8�h�^R��Aq̮�M��Q��W�J���^<eU���ʱ�i���SWbf��!��3C�+9����} �۶�@��\ �H/��~�W�����H�K�3�3z��/%�Ô.ϸ%m#2�=v��W��<RH���NT�7���3Ul��F� �A�q1J��GQ�Sd2��L�/�σ��e|P�B��G�3ɲ�����f���Wk�'N������Y�wr�>���B�|�s��ё��n��e&]�US������P����ہ4���_�\�I����3�JMJ�>�{���)���Q�l#9jz7�H���S�٬(�p.�W>L=W�Q��9B���x�8�cN�k�vhH�k<z�I�ҐN�<9J�xd����q�d���U:�ZJ/�Q���ڣt��Y�ہ�5�$�^���Z���H��L�/��en��r�j��zI;���ч(�����2�����S�m꾞�j8h�B��.w�J���4΋�#���-���q�PZI�2���$h�sy�i^������$�p��r-�I ��6��4ĩc��X͑� p;"��<%�U>�(J}5�����u&������.��4|�r���afᎿ��V%	\��3�x��Tc�-KK?�(M���ҏ��?��L%�V�0�o�ieù�g��o���ķ 87��G|��_~15g�2����6��o2���	Q�*�1}�����U���f�a��}s����TO�*G	�}w���K��wt9{!�H�CH��f���և�>v	�~������c�8������*h�����AsnB���{;L@�Y	�7��>���� I�S��[U�nvIj��w��z=�6'�(jN�����41㵼i��.�CsfZ	�Cu���!y8~M�]��/FHʹ��y��1���@�s���2�	I��
N:['�/��H��̓��Dې`�M�\sqZ��8	{��ύ�N0�Ntǔ��<���}�)�G֫����\�v�H��5$2�]
��Ɂ������P��SW�"��V3�f�:��M�V�	��fR���6��U�*_h^~�^G�@�\.���F��oA$ͲU��j��?�7��)q��pm��Sյ?V�w���)���b�[ri���0�J�O��+���3�ctl�~��,<�����_fij�h)=��q �W�۟4D��x�$�&Vz݆�-$�⮎UI��D�(��ۈ��x��7�J�7^BD i)m\�QR{�ZU)�TSF]��V�^޻-l ��b%��M=Jd'��)����bމ����M\�2;��'?���T����]�o�/�c�͎�UM�~f��Ŏ4'$`C}��_��\�/�H��=����ing�l���űO|��]����h���5��� 5rآ�;�C���:��r5*l�9dwD8�������JP����W>7� '֮�]O�EfJ ��N��8i�IV���0/�ZU͹y�:��8��ZC�͋���ҁ��:����-�(ڱ[&�4%p��D���?K�M��R��,���!�8+���_y�Bq-\����Q��~'`q�K�R~��`f$�R�U�"��g�8�Nw�=�9���S��0���̨,q50��ňn�!��ڕs��>\��zިc&kl�*�yҪjy���_�ry0&? �-r3���8�y�7_1k��ѥ��=|��_W�ڏM��ȷ��$�,]���X�sl�n��ڽ��A��"Vq:� �C"�c���b���i���4s�E�M&�>6�JI��^r{]�C���:\g��F,|D\	W�ҫ��cэβ����D�������Y�*e�&E	�P#'b�*�#�=�� ��JnO}��R(�5醘oRj�*;�8��yYI���qȈ}#���)�����fl�p�������`�ϴ�lK5e�~:C�]�>WZD!��y�\��@f������x�D�:��X!��u�\:�6T��u�~�x��_\9n�����)�Z8��iЧ�U�a�3)��N��i�lhy�\B�pؒ�	�ђIm�S |�\��q�~z>8!q�-��OV��������T��_� 15,�����ܵn�����_��ԘH�p!�u��$�,؃B]
u�)��n�I�,O���[\��?VZ�:���nr.��|��t�3^�O͢Z�A�����KO�=�#�I;F�[������7�!�����<��7@�i���Ī�)TQ9e���8�iĩ��K� �3T[G�(�,����|�	9Y,򮄆2Q�62]�Ŏ樆o�-hZBE��ֵ��vb�|a"��]��BG�q���� ���e��ե&���c���y�%_q�Q)P܇W~o<�pP��k9]�������;�E��1߿Q�u{�Xo��=�5�<����#DDR3Bi�oq�Y2 �2�Mb����| ̑�	�[m�1{e�U-�T�q�d���դ����@! uoI���R��X}�$_�������N�#�;�姊~�?��{?��f�X�i̍*�C�z6������r�t�mkO���i���%�K�`�H����ˢJe�-��!eK&�2L���u�G��ݬ��_[�]Gj�b�%C48�k��-Ϥ����};o���H�k,ȓ�ʲ�Mv�U�ݢ)U⍳;`S;�n�����$>ŴF,��>Mw�H�z�U�+�G�mj**]I�#����Rކ�h'�/q�W�#2�ߣ���!d�u�P�B�}���C��z�DS#�׾kn�uɈ��->��lem4l�F/�)#�
��8
�����y� �Hp���#/���S��Sh�ň1���\-'Յփ�$a2���H�Y�-�`�����%;��=О\u3%Y���*)�<�s)����\����z
�Hߟ������b�i��������~�d��r)�*�eTh('t�xJ��H���Ϙ�v�w��e}��.�+e�t���2�*�H�n�����R���-I�����������
�/O�$#V'�N��y͇�<~Z�_d�߅�hV�p�5���-�j$Q�Dt��.<������Q��܎dDV
���AZy��ɖ��ނ?�0����pS�W����K�&��M���&�kN/^s�;\�ĔK���"��]A0$�q0	�[0V !�!�Pb�����o��P�����Z�S�k�J��`��{dZ�]øk���rҁI)��^��,'�������N^�mX]��6���v3o�+U·5�j�G*�4��4B��9JY���U�a��xn@-*k_i������u��~���h�����v�o�r\��(��#������4@��:W����[����aHE�%��H�y8�&���xj$+;�Pc��#�k�TT{�G��T}���=�85*��߭�p7��{���B%���z�����3����J�1��I�Ǉm��K���#8`{�\z^�k��R�B�S��uR��BTmrl��aEϊ�I]F~}v���/�w�:���]��T)��@wc�[������Yf?w$�'�wNu��
�L5L�u%���-&F��cㅹhOe.?��/�<�+?ݾ�w�ʺ�1 ��S���� #���O��X������{&�Q±���s�O\�s�V����Ye ,��QC���	���?qE}���(x��<� )����{���4���9-"�^�a�@�x�\b�K�B̚���g��h�I���SVUgJж�y��D��1�L�Ţே��Q �������B��QM(��[�=�br��=#L0+O�>J�U�f��j���K�%�ňB/%��B�b����ה�I���J��;��GS����� B�z�z ��G��X/��̩w�rK(�;�9��w֫[U*@b�-!�v�4CT���DyՔ`����j��Vɼ8�O9v��!}�8O	���R�@+SI9��M�	�%Sv5�v��$@�M8�IB�>P��c`ô����k��iJ�Ykd��xA�@����ǩ�_���Q�S΀Sj#	ur|Dg���ӑ��5]ic�=r�qi���h
㣾�����i�S�C0�UՃ��^y�x��` tj{�(X54��:����A��W�e�J "3b�.��s͹Yʒ�E"�a�͹��>z}�ns���uU�1W�Pzh)���3C��,�+�_�E��*�_}��L��I���֤Q�]tED�L��;JYz��lJ0��������Kc�Z3�&c�p���~C�YP�R�{�y��Mf�m{]vI4�Kc�C�Pf���t���~=����j�\����t�+q�4U��������$�F��F�on%@1�?�OS���F����-�C����c���r��M~�)n%�Y���Z�(�HU�[�D�p�"�gU?��:��9���C
bG���
ɜ.o|��Wku}f�U����\��yi��,�O�x<����48tTd�V[ʮ�j��'q!6�\I\��K��Q����HD Ӥ<"�x��[Cֶ�IE`�x9��x�h�#�#�|.��d�X�@�[J��BfW$$����������H��#zUJtO���+*^aL�N�R+9j�[�ەm*�W�L���[
(�	R��ݕ{$H�[���6��j�����G�����I��,P@P�GX���r\{s�F���yO	_1���dkIvCNS�r�媵-�v�T��]���Gi�WQ�ϗ���?�HN����J�B�G����n�y���$v�	"���_�U��5�Szڳ4�x��'b�ay��y"7���/Z��ɜ���� ��8j�&�� �\#�/`=?�F�$����Lجe�R�����g��'QLC�� �z�4�tt0A
2[,?.�F7�SA ��ہT��jL���q�D��U�����Fe��τ��# ���p'�I5?�E�٨�����\Cq�S%p�Im��)N�pg~}��݌���N�S�"�����[�ju!U��낋��?)�ܻA��c�u�uֽ�qP� ��X6��$fش�=��#($�+��x���c!'��a6��M8�^���C1�Rn;�h�C;N�h��D��FzK&8x����{���z"h��A%���iR�{?=��1��ý� 2OR�,9j
����ɂ����N�" �e&�Yݡ)`�G"5�>�и�{e��a��m��V�'&h��yeX��i�F��;���iN
��4�]�;���X�qT�)���u�)�Ư�)q��-�����ڬP��1t1GaϦ�!ߜG5����F�ұ������_�>e9|�Ll�:�ɭ ����o���tV�9��)��h-���l�E�r�8�+O�/�^K)���1�]
�ć��r�y\*Vc>H2�A?+�MuQ��kfkl�m�Seq����ߧ�7��T .c?؅.lN����NsTSq7�?υ�&�h�[欲�ބx(G��y�!��i��
>�>XfcA��♙�����Q�ф#�z��hHv�: `:�w)�����_�9���!Ӌi6в������5K��t�$l�)�1������s4�Tқf��C��
��~���b��@Ɖv)�P}cq���hC	W�X��mR���.�ig.�#d?%(�>UE
S�92K�t	h�`���xMO��_3U���T�@@~R������E	��m�C����}�S�\>���Rт���݂h��M�c=?�Ng>o�h�サ�8܂dŁ�Zᕱ^�5�$qE�T�wmq�q���n���e�1h�[�ܼk��MXOI��A��a���[�"u�8;>d�_*����p��B�? R'�:�s9b�����~�kSOμS��(RZ�;�(�%3n��Kt������ ��Vv�4�46�H ��~q	�b��qG\~,�`m.�& �9�"k,���J�A��x�L:������t ����Q��.4z�7����%ˬ�b+��b�`m��j�!8������P����*����ҁ�@�D�J
v�l����`�R��C]�H�o�׹�i�K�	�Y���hZSɴmr�s^d_�O��Av��7�1d�}X�:7)q���~�5��_S��;6��o�{l|���_e�����鏯#~=W��.�{�iS#�*��=������;����_ΐW�v�Ã�[�D�=�b���-(�x����uz�}랸����]�{���4ޡ�^[�pZ�do�C�&���]!;��p�2j��i������h���΃.-��#���)eH#2a��՜0��}щ�V\)K�I[��>
���J	,%&���� ����g��N���]A�w��[��]4CPa���l�r�=�۾h�zrv�ͤ����l"�źU�J��8�޵���N�/��W{r�*��_�{���9���.�Dc)j�\�C� 0s�*&����-�(*��j�hQ95����P
�	�si�N�����i�G�"c�m���%����26Q��[:�'D:	�ϳ!u���̌!b��Ő�	ǅ1���q�;h�x܎�/�շM�x�_/�f���)NV��"4�29QN/V�� v��\���ϧ]�4�̕�����`���V�˂|�&�;�j�r(�#�/�]]T�\���Dc��#�x�=�S��-o�3�G��'��=�]kmy,��_-�4 ��ʘ��k�����HMVz_0�Q��w^?=�d-д9@��Zܔ��������"b��XG٥�	̰���U���v�e��KXXq�n�y9~��z���,	�W���T,��qMJ��w�ue�"�W��949��ƶ�Lq�[�:�҃�Q'1�+Җ�l���*/�L�������Ȱ�\K)KDo䙌�6�I^2�`P5�d��ۄo!%g&�M�'���i���F���\	�j�}(_�6M��	|H����_���d\5�e󌿁Bá2����&ꩲ_0oܭ�@N��;5�l9�����S0��md�;��`W�83�oL~P'���8{08��߫�0^`���QWKR��=t��G'u���㴲�
=��&���cK�h����c���v��WZ��Qw+��t��W���:���]�lHZ��Y��*�\$�c��m=ה�mo��Z@�t9��
��)b���e�0,���}	@�`l�=h
�%��1+�p΍�ȥ\�-'�;������IB94�Q������E��
��@J ��b�F�,���e|�<���L̝m�Bh��5���s?͔<�.&�3VY��b\=J�%�o�C��LoJa��:�*��m����� �����}0����|%����w]Nng�B+5Օ�w�[�f5���y�û���\�ݗV4z��!��F|>3[Ғ�D}�"��(˔�����G��t������P�9VNN�H�������+�Ȕ���da����m�W�c�We���6��A?˰�S*�q�ޘE݈>^����<�����4��� �cܩ�ؑC?�n}ǯ��?�!!?Nɒ���M$��!k�v#����gRj��d�1�r�i���
n]��!T0�T>M���`�"M�l�s"���lq*w���	���=��c�H՟� "OH}8��QӜ�r������"=jΗ�w�0�mFd�ո���|jl�d�d(��HJ�^��T{����e9��j�s.�j�#�_[U�I�4�üDb��ao|k�8����q���_��jr�9U�:��Q]�V����^N�^��iHs/�3�.��y-�!�Ζ�1����|���H�_<�&���_��˄�{ґ`jI� X�Y�.:�.���'�������M�i�����&`�4�j�`?$�{�/�GGn$�g�X���m���6=���K�<�55
D�CUz��*5-O��c�{��G�u������r$=1�����/�چ��n�� F�/��Bh��Zc�TN�Sώ�>��{�>��-�DHǹ��h��v����-���C=m*�'bR2�-��or�Ò�K�f�\0��Ol�95}�L��;���iP�4'�w�M��꧵��^���a���7��&���]W��\������3��Xzl�A~��%;zt�h%-EQ�ҍW4�u��J�����C"���jv�;��W�r���L4�o�ڑx��� �uƕ����L�u���vgHGP0{�M��߳N��U�������dЎ���mH����͊�º˕���8H���w�?!���X�(
�[�CA��2�o2h�k���ԛ/�/@-�7�{}�f��}�ߎ������VՁ��~������P�:;�=Y��~C���$��ȒZ�o�S��R�$A�����i�V��\�"p6m��\�w�D0Y�t�BZ�z$�1/�V����¼AU�*l>2�+��9t�D-�k�e^�Tζ]֡[S���\��#�@����j�_�Q�kL��
C$��oUޏ��!�<�~}l�������K�
���+��^��6�a��[�+.\�|��	v������q��b�Yn�VȒo+l���-3
��?I�\��ӼΦ�)g�f�	&�"�b�9�uF�����¿e�b�U�I�}���"ɼQ��)	_�/��cr��IH&a�H,<wx��r�MM�����[_�|_���F��k��a{�.��1u:@�t�ʐ���ê?�vY�BA��s��f��r��qZuܑ����d+E����XLM���Pg����?���$���G;��@_:��oT��e馢*=5�Ƨ����@p���p���("/ز~��z��8�.hQ7���9>�H�%�>�t���bMD�+�Fxmt�YN*o�3�tå~ {4y�E��P%�}���㰵g��׹�&��׈	��2+��K��o�9�������6����єDZT���]�7��1�����Z�۠��^�h)T�W��5����!b74�R���0��6�<n���`%}������s�K;�U��>~����SP_gD�Z�Ò��)�w&��"�K+:�sC�� )�����"t�v��gZZ�M���Ʌp���"X6�׼�9� ���JZ�6��7��)���b���ށQ-��F>���5��\n�+��A8���T~N��&ط%�z���|-�j��l\�:��@sD��O�t�-��K�ep���-�U��(�]���/祳����"H�m
0�e24�񆿲�ND�ٺ~C� ���T�w�c�П�:�D�4ؙ�i��<�[��6[vb9�%k��k��)ݓ����2w�(��M1�N3:=�MO��O�# ����P�*�С���z>����EPtZ�E,ĪY����*ؽ�n������g�:٤��.�5��c��j���E���dЮ}Q<���BD���ukġOҔ�=��V�� ��$��Yepv�L���(=�}b��&`I��ez���A�}\��|�#�|	�^�\c�ڗ�5�:WG�O;%B���"a��K�5�I'�`��*�v�k�=k�Sn�z[.B�����g�L?F�W̟�����SVi{k���*=��l�ۛ3ىJ-�U}soMn��>n�Ꮧ�,�+�Q`�_�]~p�P/'8�dS�/�O���{��������o�_<�7m�h�L�9�z��&B�b%N�-3��$�����@��p>-�7Լ�;/�q_Mlō���k/o�L�������0��p����1[�Z�6���)[�_��/`5���9q|Z?i�~I����·���b��35�[m�ƭ#sC������Bߛ�����Q9�^�b�tԣ*��\�v�o�2NI� )�|����|� +�T�P��V��p�TV�u��r����r�QdI B8!��S����t[زSΥj dF� 힏�ǹ����)*K��;�E��$I�k۶�uc��PZ���
�_�AU�2�܄�,m'�K�Y=�`���#19�ݺ|����a���(:�x�Q@�u��7�����9��4����6���9��wQs�g���v�L��Vgc�HJ�;Z�O.*%�0�kK6�$��OYQp�F��08����av߲Aj�)��vC�w�D�Q$�|x�����-_Re�Zv�Ԩw:d[�^�&0��M%.��M��Ϲ�P�mvf���<Pl)�*��s٧Ҋ��j[���x>A�31d��a:r����"�I�7h�(D�n��X�"c^�VS�z(i���.��ց)�N�ׅӝG�����N��aCj.6���A����C�u�����-�)ӈtC�iV-�_u6�n���p�nU�	aJ������#%0��tO��=�� �3�4�"E��[�+$"o�mjx�=th�9�9���M�و�[���e�ʽ�uh��k�mϮ��ʓ��owyӒ<nB��'���j6W^���|&N��:S'8y�������cP\:r�5��=����p�~Ϲ�IɻC��yr���̼A�~]�o��n^
�g�O)�m�<��Z#�΄.�,=��;!�X�x;�j����b�8$��J�=�n�6\:�������pO��+�%0�D���	;�l��Q7,�EԀ�m.�;��&^��~a������m�G�qG�t�H4���|�82KCwf��P9��|�x1�:��B���Q���iZh�^Qb�m��翫���G3�A�.�&��j��{c{{u!�J��{�Am %�V�?�z��L�n-[(���*�F1ccje3�iu�fY��;<�l�-��-*�Ł�CC����Db�Y���i6|�u����8or�
G�54�N�h����|N��5�Ź��Y3��T�\����
�P�ᄇe�1�3��]�s6���,�8�B�a�-NL�q �����@��h�e��K��3�����DE��#]�m9�ꮠyٌխ9�Lz�Pj���6�as���;���6�2G����udjB���!i�j���(i�E4X¡�l����Ġ��7{X���c�v�t$6�%�rĚ��g��e�!��� ՠQ�2���I�H���%5K��>�R}��|�w��h���lvOH,n�u*�İoܢ<��P�{59�����r�K�^XR=:S�"�Gl�:j�.����}�?cC�o�,X�����#VԸ�ŋU���L(G�DXr��ö��/k\�Ku��[�սt�~�ˢpr���:�1K���,{w����1^m��T��hH$}(�h�lb"�
����<�Ά�m��T$j��4�q�R͐"�#{u���ف%�����z~4u"�x~�O���n�<��s���-ڌ"5���Y��W�O>i2!x�= �\�F�ڊ�fc@�*R�u�� Х^�Pƽ�46F�ϛ�2�F;��QP�~O�C��k�߶�.)��<���Θ��xŎ��I�N��Q[�a�Ņ�����h?`��A��kyXP~s]�P��k|�OKx�ԃ���ŕ�On�;*���w�K!G�$n��a� o����Y�$� �I�r1�R�0��an�2M7+�Q~Nc��E�-��T��s֝��n��e��_�=�c�$�lWa*���_1qÀl��>�Mh)�M���g�q�+��o!x?���X�@t3��C�JLHd��}��T�v������hb����X��+*��'��+��?)>m���ⲃ�����Vb~�M��PSB<E�:��GMk�2�j����g��*�b��p��<�%���d"e3�t~��_?W��n��N�y'I��u�*���S/R��;D��k���ټh��_A�Oηx쪷�y>�#|�A�з���eCB�Á���O]2�|�ɰ�WH>��Xh^N�7A���MTyםVT�J����(�+��ӥ8Ł���.�6�������)z�a�=�,�0+6�	{��@n�q�Y��":������g�g�dP�@qt�q �oE~xڑ��7 �`]q0Q�Й��t[�X�p|�<y͋�uI�S	��W$�Fj.����"������A/���y�2V%`�ʋiۢ5�-�竤�nL�l��D$��T�>��V`�����`�aa�#����T���6�ɲ�J�]�d+)k9S]��^j:w�;4�}���O�ZƁ���tH�6�T��O��{�WA۬oW�e�A��5��9m����Nœ0����L@6{�	K�G��1�L�c-�����]�DNQd���8�w-,���E"3���^/@��8�%g���Q����/p���=МAu�H��<N"�?xHmm|�t>����0�&}2}�-�5�,�d�l�e�?�I޲�p��/'��VE�����eW���Ϗ,�� H�n=Wl`0F�G琳�5^fZ�m<��$�������r�t߆��A���Md�X5�p����4�
TܼyS�x@y�'�X8F�X�|!=��v�H�2lR��?�?l����H�������{@�̭%4j�4������9��,+Pw*�˯
U8O,�ټx�
"kS�5��%�u�y*h�/�YV��(�_>��3Į�}Cq> ��=�p/�E���]�3�l�z��b�̿S�\���ҫq	!rAG�BЌ�:�P�UP�q%���m]�8�����݌3wũ�>d]7/գ�{f%�Qҩ�)	���Y���'h��	f��
���Ǟ � �ҩ����m��8����l���O!�RT-R"����]0��%]|;�˜b�z�YYB�70d��!�e��/݇��u�V�[5v�����WT�C��k�T�V���S��Uv��@��j�Fξ�Sd�7���cg���O�ڄ�q�z�z��2.]�_��Z��,d^�=;K�\�,��үI����&�\�#*��̝.Ub|=]��*KU'C���n�>h��v%�2�	�R)9d.w�C����s4L�	E��(�֔P�˿�/=r���C�m��˒r��vү��A�~ck|���$��`�������ž��.�G3<�A�u�����{�x��_��IpE{�U�a���	��[_��|Ȁ4N�.у�W)hJ��@*��]ҙ.��/	/bD�P`ԕ:6Cx��#�Z��L�RE�lJ�#�ɾ��.��P�e���e��/.a�0������ ��=G�>���N��	3���E�˘H��em���wѱf�U9�XO/C,�� Ed�r
LPb\٢q��ضM�xx���dfC��CqG,P�z.��ج*����k��tʤ ,��Js����x��J�qU��C.Z|�+��Ɩ��t�\@8��=�Bk�3��8Z?��O�˦ԡ+�C>N�\FĪ@�t�x�I��LhS&�]���d�S_�B<Y�b�V��B]�:���`7�t-DiYX3r�#�e���g�8P�^�Jq@�C$�E�`��@�O�P��,_�T[30�jE��Dp��C�Rq��]o����J��d|ڪn�/W����܁tsʸ�l�k"��ɔR���vB,��2�����Ȣ�Gum+P�{��i_�L\Hh�t�F?�s'����&������3b�s��;���.N��&p|zJ���8��\�~9S��VY2��ol�.�����/��y�=��o�g���FfU�Q�T��Jw���pы��8%�e���%�i�8�$��w.�7ƃ�j�+#ɒbs�_���f'��j�?b�����ک!~̻��{����Ac��3�E�&�;Ǝ�BԎ>!ޛ���eUI��Nx�1�>ԃ{��S�Qf�xv��+����}�_!�dr�d��&&(�P�Rz$��������a6��"Fttx�;U��axB
�������U�3���b_.��)�F���<��wh)	!��&���,Ӌ��HLW�$����&Ȕ���y~T��]x���l4�Q��t��%|���{�
�Թ�(�x�i>��R����hlF���e>��\F�DVڈ�]���� "�jI�����6��J��	���^��1Z�v=@J
��7�/�[��� �>���	�a��8�^\���&�u�gb*�x�Kj��f!����G�
4͌#�T�sqWmZ��H= �!��fFq�<��Ҕ��v��T��J�,�1��_�P�-�(WnZ���UL�U�9�mU%P'#�>��C;���\��n���ߺJ���/ɫ�ݒs,����q�y�[�O��/�m�L�gzʮ.�B������� �F���!��~v���^�vq ����5��|����}f��O�m�~		�2*�8 F����?FY^�s����Ҁg���(a�J��������Y�;�w	��0��"�Qﴂ��zz�	���W�˄dt$��ۼ�"`���0�����v�v�=~0�xÇ��AL���ʃb|�"��Ydz�����������Dx0p��i4tH�΍�O9`C�(C����n�5�6}��e;��d.�C���zK���y���)Z[�}����3Zv0۞�k��;�����o��ȥL�֪!���5�b?�(|;/<������x�`�nv�u"!o	��O��Lڅ�%2^�$(@H*�V[΃�}�u��;�Ь�(tg��(Վ�u�g�I����ƙ/>��a2��7�0���@�x)?����Qs[��.�VT��u��Ȥ�E����]�d�-&J^�.�+�m Vk�ԅe�2S���j�B<>y�����D{�"����3�[*�s����ɫ@x��m�����%�������<1�<�.p���}_IFA��]��<&�"�(}�������U:���O��%y!&n�;���- }����g��$���8�lW���H�.��w�	�8�vؽ�&,�'�l��ƚQGd����V�	���縠��Z�?�h��!�� �=_��B��¢�q��#-��--ko&���8RxɧL=�7�ݺ��I��	��W�����A�ov�z�qs][*ಝǪ�����[����5�q���-�nF#�Q��VZ�z���-?"[�~� �u��H������4��E�z��ǧ�C3�ǀ��u� I�l��'����u�ݶs��Y��Ǩ�plhģ���{n�����tݛ�;����v��7��50�x�!j��$3[7�a���y�"���#���O�^r⇬����1k���FQ>8���n�h ��v36�ue�W!��[�a���[���[�����3�#,?�u[���>*b���E�8�ÁOR��ٓ���%��n�J�g3J����sŶ��	8fxF��`���b[�Kw`q��~ּ���U�l�3k�.K:2��1�]�۞�z�6��.�CEX�ʤ��O�,��S�������7䔎�?�p�l|G�4#���+�~���q�<�3J�2�v�g�Ѓ�o �F��j��fs$.�^�!�k���I�"�y������OU��g�Oߏq�װ�P 
�#�[.tп�x}C�(wݯ=�Zs)�],Wd�S����y�׻j$R����G��{A	ʊ4κa6��+߱���Ȳ0�5LwUA1��Jx���?��"��m*�tl�Z�:Z;�gVl��Z������-_���;U���z�]��mus���u����$YvȒp�������4~�2�k�c�Y�>��y��+��( L[ȻmG���a�>0mM!!��k��Lװ�F���^���6>�4�h�oG��U�>��gV�eD�y�,%pm܈���D�����k����?���>��&V뉕G��C?7�`o��n|]���N�T![�Te0ק&��ǍA?3�x��+���8�����V����Q�<X4�ࢿ�%���y�d��f�l]�1��C�}��7D�3A�L�η�fuMFp]��,�E4�`Za��:4}BR{�8���$R[���4�S��=�y��x��4g���u���J,�U��n1��?�m����aS���x�3�@պ��|C���2�r�O�r�ĒA�<�o`l�6�e��-QI���|?[��[�c��S�Y:a�������U������c)����lDr���Or� �o��*��,�J�>��\�mU�[BCm�9X���HX	�&;����%z�)<�ȟ�xh���|qN���/5��/�"�a��RghPbǼ��f��J�HT#�|-��&z�ʅ<�9��Z��x�\_5)�$������s'ʑG?����|��9�uR��O;��&��?4C��\mU2'�a��:���O�zcN��:�?fj����.Q�p%`d��z�-��	�7P���vz�R�H*�a�vE<��hl�_$��<�0������O��q���j6��j��]��艰�Fk�C�l+K���K�V�wO��d[%�d��%#��k��{�9Ht%JQ��!��kۣ�ܵ,� 8�L�h$Ǖ�.���(���Y�$����ې�^��O}n*?���]�G�m�$�WK��<b�36�����vLf���%MT>�s!��9ڷ�9\7�u�1{�gA��:J�����Vv!�����#
+�:�!�M��x�auCnKS�=x���b��tҧB��Y�F�z�sf�-bb��Z-�����Y-�^D�oR-�����s����������9�'h�7A\�a���n���� �]�\^ɯWL�rZ+Yn�\S#�����2� � �]a��)o�j�������r�������&<�}��O�=I�3��u�Ca�
�q�y�v�.�֍,5i:��b�Sd�e�'��Vɧ�&  �[DR#���9�@�[[fRǳ� v������ʙ/@�rOX�/ɟ�~�<p�K��KCOr=�t���il��<�I�97 `� ��'3BI������0��u@O����	w
��t����s��_�z�Wz�A�\�	�$��<���O �1.s��Q>`�q?�ɧ��-������^_�怗���b8b�rO��j�m~ڙ�>6e��J���X�{U�b�#tFKp2;�@+����J���F>�ܘ��+O���	k��s�>����ej�^e,O��?�-������*	Q��{��-�P�۱�~
MI�ef@]�(W��H��c�-z��i�ot�l.�^�=xV���@|��H�;�,�gd��}�#J����B��c=���QLĭ-J�3�VO\f)�q��̴c�l�o7pp��������p�E!�D9�ۑ*殜p{�!Aߡ��o,��R��ͧ�e���w��$���d�*u�2J:�7lz(�����BH�sԙ��.�*�s��7��8�$�<$#X�9���)�N���/n˓}f�Pv�~S���E.53���r&�(i&(%ؖ�g�b�` �3�kTu%4\�W.�$��U"F�lB_��Q�I�
>R�k3� ������!^�zN��(��SeV�mJ���Ӹ�I09U�KN�B�m3�SW	�"=K���Kŵ}�M��x�e�̟YĖ�ެ�u� �ۇ7���,v���	�c�� �,> �ɽBu�����}l�����Ԩ�6{��Ap,�]1���qW/#�Ʉ�/�����|nZi���FwRNn�|=�͌z�S��i��g�ΰ���$[����g�hf�R�=�F8�vb�S~�a�)����#�s�D�����<�����ő�d�>��*7G�HP?Ɍ��ɜ���k�^��d-�d��$Q7�Jꀖ���!V����o�H��
��	�T�aH��T�P���Z�)Us�8�����$r�V/��/�꾙xZ:�{&H1ʖ?p���Uh���9B�UJ�pF�����ԹD��S��SR��x��I�}3	~�p��7�k��n�r��%7�������'���Gukk���tҨw`�
�Ak��Q��I+�҄�kZ�������g�������C�Y��ΰW�7��/lf���W.��i&h0��<�q!F���H��u.-U����ms�=�+�cb��<�f��_�̤q���I�����Kʠ����r��N|b��d~�Q�~$�)�[���AD�tUY�iA���!��wW+*&[]�%�o��}�
�2�ݢ�d��;��b5�Tp0$��C_sD�&}�a���M}�R�:�9�"Nq�ī�d#�jM|��ۋ������=�,��Jn��,�G�K[��-1���&�h�����eU
3�&����Ԫ ��~�)vz��5<W�jh�O�׿
Ӂ�,��&/���k,92r�V�&�ψh�20� K���6�.�A�,��;N������mU�9N�X������� �g��Qf����Q���<Q>/��yc�8O�b7��:�0͉5�߃2j8L��ʕ�?�j G��/���Ep��NWH��`��.޲xO��P�+���R|]T�t�p\�5&�]�-Ц�,	z��)��N���F.�c�t�CB6����t�-��r2J\
�c0��r*���Q#�e�M[(�5�6��^�Oh��?��"�u��̈́�S�4����r{h>y*��V��L�=p��oa��ݽ���4�4�jOD�mR�5Pi��f�!S␿z�6���iL��-��<�+����5��J��~���a����MC�~~���Hü���S�E#\1���S!8�S׻ %%d3���o\�k߁�`rq2�s��v��O��90��:��ww+��a�+���cd6e��^�F�2t9%����~����2߭��f�,�*z�!��%�>�
z^�I|��!,c	�?6Jpt�~�F��|����������V�p��k.9���(#?NÀ��~7�=�&��܌�^KU�vN�pz�]�3�l꤅+'e�q�Y{�<KO�\���4���2�?4���TO1]�Uo�������[J�M�o�� ˗1�y�����b%X�����&p�lYb�h6KCp��� �U~�d��IO\p�-C���A�T(3�H��i@==�.)��tN
�_�N�-�܄�_�4�g���7�-�(���5ζ�.w��:�v�p������^*p@W�	�i�)TY��"xE�څm4�z��-N��x�J��:#��8�Z��s6�ȝ��X_���H$�E�U��o�h��bd���S���A�� ���h�qP��	P`F��Y+�h0N }�lYj!�f| i�|����يL�J���rS��ڧ�\���8���=DZ�oӫ���z���S���vA�Uظwvg�]I � ��m�뢏,b��
M���Y��ҊOS.�#0�-N�*<��k���:�G��B��1��a�Q�i��ܹ�acp{XT�v�H��S��oT�֡1�R/���G��P���N~�׺&F^���|ב%�|�v����)$��L�!��I��o�Q��~OJ�I��b�-�G������\)�g��Tv3��-�:�Y��f���OEO�.#kqG���J�����B&�drMW���KD��?Z��:�{��\���^��~�I�s�JFT<�uF�Ș[�� �`��x{�۸R�R� Kur�#
E�kh*�+Gs��k�z��b�����V�-(j��:�gP=���+�E� �Ȣ�g�8X?�7�Lg��V7HA��(T��c��/�>&d,�_�6�fp�{(-�ݵ`��h��'�)!\���$��*�� W��O��pW:$ ?_�tKNb7ⷕ��U�0u�?��M`���{���[����E�B�ϣ�Єd�Of~������*X��3�A�`C��� �XZM�]R��{o|*����T0��o��GO��nl	N{۲�9��*s 8U�O�O�C�Vuw��p�Ǟfy#2�g�Z�xE��bX��Q�$Gz����"����B��3��V?��+I��3��b6L�U����o1G�D�`���k�/Y��cv萟O�Ϻ�|rr�ޕ��P�9q-�X{e�6t��@O�;'��)܊�l�t��Bݖ{��7K�j�������w���]�@��]B�M
�P<I�6�Qr����~Vc��x䦯�F�< ,�3�<G� ���0!�8mf�'2�ܤ�r�M�u���o_i;�j���~�JBG]��`FF��GA�d�+d|�>l���%�Ie�h���U��(V�Hm���J1���ړA�n]��
��7
�n�̱��W�mz�oY�n�ʬ�ej1K=�0E��������0$�x�id
y���<�Yxި���	��(�O�ڰWTq��+�"e�;G}m����/� 1�̡�L��%S���4�k6�㸘>��	k-b�u�oPoxo�
Y Ɉto�˨�D���Ү�w<���u�.�'X
5�t�ߤ�8��gr��F�/���T�m�:���N�K��N�!�;hD�Vlqz�I�ޯ�L{��O�G/�F�.���iL双���.Vc�� ��5V}W_����ppnc���eGM�H��grkD�Օ�H=Z�x�3|ۻ&|�	pK�5~]�����周�s������h�yT�q�S
��xR@� #�hm)�Qew�*r3��l!<5j���B�)�GDL�*�i^�gF��4�o��å�s��Y��~��6	��@�F!2
�����KR�I�H���P'"zd�M4ՠ�|{�NRb���-F�
Kq��>�Լv�h
����:�Y����}m�B���	������r�`�(M�'����*G|F��Ru���+8VEUd�9�&S�A���z�d� ��Qٯcn~>�gs�צ"��܅�	��m�����l,z�\=X�VQ��BhyR\äjs�E/��u�T�j��Տ�
��m0FV�Y	�F�i�Z��f�X%RՄ��H��	���e�Oa�ɀ��<�{&ó�Q���3�A@R�i���k���o�,b��U�)����v�̀���Z���S2��][�Eܕ�7�Ly�X�5!Ƀ���&Qk�<-�[�5��S���D�g�"���:�'��=��j�ڙ��罃;z���E4+';�D8d�F5 eBJ���,S�R8�w �e���4�J]䝸C������	�pT�y�%��e2n��x��i4�H���~ӱ�|؏�+I��{�?�����V��1����]����I�t���VJ9��K���lVr�7�A�/� k�=���	=��
��i��9GO�JoI'(WZR�#���r�/�+6����c-y��7�~Q'��+r���=>.�=��.��#̞a��չ�����U�:�Hg�Q�$����;����S�����{��*j�%P��?�X1�Hi"�б镙��\���9G�8�
s :u�y�X��=%�8�sw���%
��m��&�5G�>\#1�J'�"]�j��L��˸Q�.Z��!�l!�����k�F���O�f��c)(m���>���m��p�l�w��-�9�(���;��+ ���(_�F��������[�M�=����<��Mp�G�̏N}�[n�?Z3R��g�����.���P��2�'���3�f,
Ż�؀�	F��v[�`��%�K��@,����~��q(#�������Ǆ��;�Z���A9-��m��5�e�,_���w*$����w��W$�l��7x��Y�P�|���(�(j�����т4S����4�P-!�Wh�����Pl�H�ܔݛ�r��q�@? p�ze��i��m��/NUF��}����֭O5��\/Gi��O"�n��X�;��e�gޕ��t�!�$�Ǌ��;��gq��5u��($���O��rCe�^4�h��� �4�,V(O}ߡ������.����7J5<[�Y�]p�k�͡�W5~�{Ј��a�0��C�=yN�~�L�S�'i�P�)�(T��1�RQ�	��xp,���y	/ ��x5A�{��ׯ�(���Tԑ�\�,;)�+W:��� [uV��H>�,���uࢬ�Cr#�
e��E�ID�Ͱ������S��{z�r��>:XxE��5V�u���\�W�4GQ(]�E�Y��W��xt��4v����$��}���r$���>��q��!������&�5�� _�=:�����'pu������ ,Ǚ�f�z�"�kޠpc�&lw��ڪ�8rov	c��^�͜�1�E�ߢg�]T�R���f��DFGMn����1�cT�z�}����0F��#}go�O,B�M��}��m��J0����A���f!��6$S\Y��G��hp�<)��;2� "(EU��0oG�oUӣţ�bŦ��N����G�,)LG\d�&x�Ҟ�޶��<<(��>ϟJ<a�$�+3�Oi�n	�r��..��쯩FA,:��r�E�k\�HK�<t�K������W�G�o�[H���)P�W>�c�C��Me.!>s�S0
�O	��p�]��`@�B�Ѩ���W2�`���'�27O,Di�HG(� .���"��,�Euh�����;c��l]���w�����	�� -Aɢ%H-~�	���I�CXN�.����9�2��焿���5}�Ͳt�:�KHء�W]	)d��x�a���G�]���˾@��[�HB���+�ډ�Li��'�( �������wKWʡ� ��}�N�Zt���J2��'����qzk�0�"�)i�ZwmԆ�Y�Z����R�)B�?���:�ʫ��?�jy@��
�V�e�,�d��{�~�ʋz�����1,�{'~+���S2z)5�i���ko4�ya����mD,˖À"��/�P:���Wg�1�v4A��Ti#+�Cr:�tʢ��� ��>��v�	��l*s�qcr֦s32Ƞ��P�����N�c�L��7l𜱸��Yݻ�|7~�5�˞�H9wig��R�o��*�AѠQ;w7�=�L|�g#K�K�9Q���1MNR(�d�s�^G���O3"�;߂�J&0a�o�J��:�S���ڠU��w>�e8#�Y@��)�f\�ֆ5W&�}�J6�O�f������i&����CXV6�<x5��5<E,����,Pg�-�r��h����q��g;Ѹ��O�n�y�ʄ��B���׹p��R���d4�cM�7|nk��8{��<��ʥU��۝m�0���:�x�ǹeo��?3�?�5��ϝˣW�f/�H��î���{
�O1`�I�:s��A�9mJ/����"�쪭pl���g� �lO�m�T]Έ�9���I�Kr2�͈]�)h_����&V'nbK��[�K=���}d\r�[��6b*㴔�,b8��14u�5�Ў�ֿ��AhX�f�W<Ji��k� Bu~��P�-�6�9��\XH��~<T��q����Bj}���I����H���J��gД�kB�a��:r��`�9[?È��v�����h���:}Wu�R�2'�}R�z{}��L��{bh/�@%�wB����B��ˋ?B�9,{]���ι�}�
���0�C�<��o`�}?�xK�a&�"�	�s��47ؾ���T��E���� R%� ��ˁ:ށd�v��S@7M�f�%t�C�|���lqo5��BԚ�HM��*�dg��y��QHxZ[d�3�R�:(���j0Y�^j����V@<�m�4�4�7P�i�Hb���&�:4��5�ԥ��.h����Ϻ3�Yii�|^�������F㚆*���?s��ۄ�9���4��;�$wOe�?<���y�+���ǒ��S�j��e5���^��U�`0�kTU��M	������ b�w3-t����0D+y.t��*vϥ���R��f62�5p�f��}s�x�y�V|�*`�:�SK͜�V|n���d��Nf!W�E`/��<x�w�S#J̮����Q�9�4Hg���Y� [B�ꌬM�( (ENkOݣR}��:
��fc����D�ݠ�-$_�jMӦ�Sʿ�Q�P߼�
p��
�uN�����gZ�Y���u��{#��j�������
��Y�J&(�|�n��� �EV�m��辡�B��S�dG+ޣx�5������J�� �fa1�
b��T۰P�ʯ��mNP�TRt�z$�l�i;'⋪�Ȇf��S�g���������
3_�*��WNWY��	:L�h#|9Xٖ�e�2�H��b=�0Y�A���@�<<l�yw�ّBp���3k�"����vg��|�dE���FֱƠ=��̶3��w�����S�^0�X��X��V��7���N^D����]���涼�i��Dze�#N�'\Eq-���{H&rV;�d�29��W�.E �_+��^��mj��H6y�;엲к���.��$�`2�Ɉl�%��e��Ԗ��]K0 WU��]Lu�Z=�/8!KVţI{�� ���_A%�)�@
�:��~���C�z"����b_����κ:5B���S���~9f*����
{K/��X�iW:v�k��]�@�	�1�>�����Tצ�62�7N���ypjLu�,��p*�ѱ.x����N��Dǵ1s0�=:��Ƈ`fq�sva���RW�_ ��(�����.��<)��&.��l�>�V���'qp_���XcF����rK�f��~�q]\r\ih����=G��;t�T�c��H&����o�fLJ�
�1Da����в�+�+�����|�7�p@�'�~� �U#	��>��=c�i<N��Ԓ�4*f�� uXAP�4z�l'��=*�׳�l�Z񦫊�Jws����݋����yRKLR���ڠ�}yu����%�T�Q�(n[J��;�u���~�~���U)3�hQ(U��-�q�T�ݝ��%�d�UF5Z�^.t�9+��n{Ǡ�f�XM��1�=���ۀr���Lq{����.]��7���D���<�T � �=
U٘�s��A�L��"2eHx�n|��c~!z�f��NG�6Ȱ�A:Йv	�g�zW�~1�.-dE��'6�P�]��w���"-Ys��T�"w�e=p�o^$�2��{,׎@��͠PNf�,�'?i�|���b�Jb�����-W
�+\U���AT/E8\z�%� ��%&�4��ٴ%�ԙ��-�hY�]���BMc��Y~��d)B��WsZi��A�
��FƧ�`��狾��Q<�(S�RP�S`K���NׅI� �p{��A�)|�"2��m�лRW�o�n̼W�l���}�lG�i��Æ����=L6H��@�3s�ʓ���N��q�X@���_6Gg���Rԍ�|��`�S�V^a����RY'-��:8���S1qs���xs@@��V�LZP��:��pJ�엔�BVTMU�o2&%c����Ƞ���(ްs�B��Y�Fj���5hm�d�%=�Y�%��7�"0��&~�BSu��;a��p��BRV6�Gw����+�|ظ \۫�C�q�z�ԇ요��Z�
D��x��<5�GY�lT��G���\�vNb����g[OoH�	ɚ�Ht�l>H�vggp�� ��=Lo�������^�$���Ԧ�ٱ�V�2�v��|��?������J�̪�%J�5!��ǭhW6K�������d�s�an��g�s���^���ȽW�=uU�	�����%8G���~94��G���Z	mTx�U`�B%˲ok��c^�k�]��&݃�G��<W���'�Z�,�Qfm��o�Ga�?x�cߓ�"Yo�S�g+����bT��t��fɈa���W 1
"��**�ɣ(} �#�9�\�QSY����RYo�_��cF�K.0e��x���`Y��@ԇ����p�Dа����>#sL(�}���c"�I�4;�@s �o��Yd�v��� v���"6��h��m�"�2,[��J�c3ߚ����<��~�eG��;DX+T1 ��V���N}?�&Љ�$�O�P��=�?���U馋8��Ϸ��^+0�(b�i�Ǭ{�+�:�$:+�b��-�q����{�Ӎ��y���kal#�p������D|�ᄆ'��s������QJ�ש�~@;6
��s�l ������e���og�~��)O�q � PPl@����Bò�j���fʱ;�����P'��^v��/��ܫ��>�h�S'B�����
�V��ʀ�<N�J[$�_4��O��$'X$����u���!�U"V�MkKH����S��k&gmC�Cy��_�-�`�:J��Np���}�p�ہV��읮s$G*�-���z�{�DvKNɡW�<�!'c�������X�䪣��[-�-��OP��|���_"����ӭo��ƋŽ%���V��Y�d��8�2
�Ur
�wb�^��aŬ|�P���>���{Y����`��.��>�Q}�xH_�0�1��$���k�גy�D��Bw \��F t��&=�#B���-�dB�^�A�aq��������S��*jU���k�����:V���_�s3]P�ʼ_�K�O�3��%?��L�TZ�ȍJ���n_�a���Nk9�甸}�+&�V���#PF�"ؗ�2�0��r�o���d�mZ^{E�O�J�#+�%�_A�R��B��4�1]���<[��Yɀ�ЕFE�G�U��������ZՁ�C�z��u�`ջoH���>��/�l�Jٿ�=h�ó���F1�j�?Uϭv��]q�M������U�;�H�a����E�`��JK�������\�,�M�����̤�&fXOOT�M��u���3�DQ�"�Z>Y�{���u�.]��Ǟ���������?�|U+k�lF���0i:E��f�����
�X��F�`��Qev�Q����Mc��Gv�ο�V��W!W�'� ���Je��[d��Ç쿎�����p���#/�Ï�SF�O�@�-~��D_��5W/�	���SgT���.�R��.U�J$�eTJ�0Y�4p�����L�5�v�J�n�8�����f�x�<���8e~����j@Y?Jl��&��
$�XБHk�zU�����7�=ꏫ�(���}��R]%&��Ȧi*PG�|�����t�Pl~4��<��ņU �������r=5m;��X ����Q](4�)3q����a'�4�ZC�ZZ׸���G�y���֫<s"6��J�&�Ţ�^��`'&�r�iK�>o�`���m����?�7����p�h�
�d7�l"7ռ��p6~�>�0��u�Kc|��M�BCO���>_����}]�,�ꊾ;A�̪�g�ܠ:څ6�;Bm��SW	�~#�Y�O#�q���,E��R ~s룊��=�R���[jAH(F�^;55�4\�L��?D�8�'�� L���X� ��3��w~����8�C_�0[�%>�vb~��Z�
3؋�[�5*��$��
�a�_ ��t� X�#2 ��Lm~n���d�;8O{:<#XYFQ���켪-E�����~��g��tn��OۅW�fF�_K�ή�/��b�zɧ	d�bkA�#������8����9�8s %�B�
��)q�����8 �Z�����am�_��m�Tq�a�]Ű����x��Ⓤ�y�>�޳�����m��G�� �n��r�u}��dkƓ
�q��
�vP�ԏiK�A�0]I�籦k��o�O��RCIi��h@���ԯJ���]J<��C�4](	�!��ѻg��D��!.�����u���X"������H������S�g������`;�z@3Xl^�(`򪲧O���.�O��
�:dH�,��ۖl~�Os�E�RZ��l��)�;�Ŷz�`�0۔t��z%�0�Ҹz�!�ǟocȍ��O���m<॑Xc���D���%���XX�ύE�S�2V�K@�$�!�o����qEr�/F���l�� �9���P��y�@�I	��	���;<E��&�
)�����h���\�F�H{ET1� U�+����5\>FiA����#�;��̃�XK��z�����l�1 ����>�`Z��Bʯ���q�f/[���O�4*�D�"Z�]R ײ����2g���o/լ�;�K�U���YjG�.��bp������bܱ��L�\�o�1�-.���Q���,;��#��_�'7c�Y�HXC����Nu2�����o� ���t�rj��w����;��u�#sVa��ρߥ���7Q�f7ظ΂���X�?�V]��ASv��B+���u��c��@�5�b�\h�WĀ��!g����G{�V�O�f��
�'(\bo2|�4ӈ��xS��<�x:�\�M��I'Ye֢@�D��N����G+3��a׊ O��9��tth��7�4N'	g�"�eqqt~&�qm�өQ��,5kV��(|�hiI�&�(�ZT��`���\D��O�09�0��2�'�7ڪ��OᣀG\�Յ�#��Q�0��҆O�J�rs��6����� % ��r�9��M!ݡ�R
�^e%]�))��{�6u���cF�A��8k�}]� �M	�,s*�z"����PE}��~�2YZ}��[+�{@�R��T�3���N���:���("qn7�'�|�p���)`�."}�Ό|�H@ٳ�6s�p�	�,���O��M#�6$;�zwkă�P�\(Av@�Y��N���"C�~�;Q6LN�	Lb�|x��Z�+�|��W���[A�ȇ���G�fG��1�x�l�uVΒ��<�#$3^�z̢��ȴ�
�z=̄K3�=�xi���)��;f9=(�@Qyj�]R��O�n�Qm����F�����t�z�!2��z&�-ʋ��j���7?�>f'WL���a�b�� ��Q]c�D#ÿ��h���J5e�����3öc��g�y��s�$�*��w�Ս��#*1[��@�E��Ա�_m� 8�vN8����5Վ^�U���;���e�fA�$2Mf�:=I�'�����诹��dЬ.l�k,O�Sù�a���2��9�?�>v1n���9�d�
�M$�x����$�F��ˍ�g�n�m�p�
R���^�l����j�p�^�$�_l�u�\h�[��h�d��z��ʚ�T�\���쁚6N���'d� �"c�w�њ~�a��4$�/SS]܎?~w�	;�0�`�-?�ϟ�)���|�@9��Sd���S:�cB���<�����V<������$$߹P�b�{N�Rߵe�r�.�!>:�!�����:I+?]�n�q�G�Q�:	�<p�k-��9�\�����U�PZ�6��a�$<Ǘu��Ώ<�F�8���:K���K�Q[�H� ���� ��F�_��N=^I��pm��ӝ׿�O�b�, ����&��	չA^�(K��&���*�i[���"�E�S���,������r=��}j9�0���zA����Ǚ��I�
-I*:U.5L�b:����b��)*��&�e�����Qܹ�$��Y��Z�&��]���p�y��f	����1]ײ� �78eo&|ӧ��6��]�����3y5�ˎFj��{�"o8�"�[fheMC�!�Ԇ���qT�P�>�=�~5!7�]^z�N2����P����Ĳj�pٽIޙ��6# ��~z��.E}��/B�߯��sAu#����(�qWN_�V�S*� >!����e�$���N!��i�Ӂ��JD�}�ω2�R�[�U��fJ*^H�$�ynԹ;�F����kJ�]��\�}O�ݵ��as�xɅuZ�0o!ѿ�8����Z(�Y���!!M�R+٠6	�XC�T"��{Q>3!X]��J���]0av���4�ZK�M�FL�3��o���$�F[}�E��pb�p�Q�GAh��P;�.���je Ʋ���G�RXo �X��������A����W�,Cu5�t��S��(#��E�_:3�w��4� :ƞ��J�MaGH�q^{YNꆰ'�P�0�F�<�~S�w;\��?H u�$nJ$�Y��`�pJ.�]�
g���E��b��t��rz3l�L|�"]��J�XX��lQ��܄-u7Ӝxv����Gy�A��w��S���dI�%��t���3~���fL���Y�=�Vdt��9l-0-�7�#�����#|�!ĵ��N�S�4=��%����V(en�����wxj��9���:��URV��=}$c*���ɫ剞f��1�$z˶d���eꚇ�W�WhձJ[#���n�ݹ��;P	8�����$��˘�M!����;�޿U> �/�5��)@�e�l�hI7~���lqon�	�m���|� ��h���=a�t6��e~xY��ؾ�su}]�����˙�/�x�d���p���gs��^]O���.��R�]se>�e	�����dQ�"�YSE�	6CXb����w�Zt�� #��l:D
�G����N	���	TU|JY\=f�T��&�&�����h�j�7�ճ���~;��X�h���ܪh����_�����J����l���EЄƈʚ,�V���(�~_UM���3ܸ2��n���|!֟��9��]c�>#�n�p
����Wj r��$*�F���^�I��jy�����y������ ?���wyb�*�����Ѯ�%��0s����#���U5�~xmy�u���?c��	���t:f�i���Þ�8�0�5���8�a�P`�qz���4��	J����2\�d�oi��#�WnQ�}'��V�)�]���g��Z�'�`��㖨3=�A�q���&3�s݀�a�pw(1p�*t����4d'�� ?�b��p�o� _WPS��E�+;��'nxx{�1zL?�z��ᗦb��!��A����f�d��oСE����_$��':��yk��	#b�Q=�����ip�o{��c�p��[J�4��Li8�Q��?����+>pto�b�4�W� l��\��� �� �O�_>����G"z��ƙ�{�6����2�94�Ј�3t��k�L�Q���&��k�ʄ��;���}#K�!1Ө��5�eX�'N�s@�1�-5f���d��y��_����OA��8�OH㚢�
E�'�+l(i�֕�6��_��,�RB׼��h�F0��L\
՝=�k�|Q��Tt�;��8�]�	���?�8?	�� �8d(�	:�� ����Ԏ�z�k��M_w�N=GSʰD��<8z"s�̀d��R>�*��9���^�����A4NB�|�Ҩ6؄�ӽ2����E����=Y�QҪ�ܱa��z�������
L5ICi�=E�#��2~S�k�6=sځVd
��;�c�|���Tb�"a׊��\��?�]�w����`�XZ0��e�\[]/�y&����_��E��El@�q>Z���_3�.x��w��B�H�O���e�!�^V5Ā"|y��7�(y����g��g(w,�h��CR�5�Ml��+���<MH�E�LCu��T~N���A��ShZ�#���ݯ�`5��v���G>�_��@ϡ\����k�)'��e��#��)��l��@��_d)�&(4���5����OC���4�S~���$�؋%�w��ͼY^�{� `�����c���Y�;�2�ǼV@g�w�}
2x�w�[�����j��o^���6�#K#���'`���?���-���i�ۋ1:Y�B{����w$J�x�|P�^�.������Սhp:,:#"�@(� �#)(S�9 ��	�>Rj���DC��7-|F���T�-JH�9S`��w�s�ne�>y�ӗ*<ˉ@I�[�?Θ�a�I?�y'���I�x�2���p<��+�+C������z�SZ;`�q�t:2�lg��g� Ƿ�ð�%�!;��3�f�}ׂ���s�ペ���{C�*/`|i��Ul?X>s��9�
���ώI&�!\��zA��G��m��\pS}gW��6�-%,9�m�l6��1�M�ʶȧ|�/��0�cU:t�,=˓6ahMQ#2*z��������68�_���B�� �|Ě�Mx����Q��K�2q����m���.�g��@�KAq��#��jgE��M`�y�İC�^ܠ,D��`�ֲΛ�0��a60���[�f`�I�?M��ϋ'������ٽ� yc�_I�WpZt��q�������۶qWJ�.O:��Ȟ��{�i�6�G���T9�5��2��q����?:|��6@%���C�ӣn�7����Ĳy��2v�ɳ�i�H��9eX����W��J���_��'L�rX�r)�#�g*t#�eOʹ1ւ�b[������=OÒO�:�5L���zѠ��K ��O�6f�4Y*�h�2�(��6ĥL�_�}����������,��C"�S/�f�uҴQ��@An�)^w|�=W�C=�=E�ߥ�u��7Џ9Q�Lԉ�=0��%�c8U�Q
bIr�����Q�1N��Q�����I�������Ǔ�=�P���M5���V^j'o�[�]�$�eA1	��b�C��W��� ��ϖ��Tq�A�J��|�g����f�7��[h#,��DwN�9��5�Ŏ]�R7x�h� �Gh�&�n��Cf��]��!�������%x���b/��NK̴�*���BV������jj٬�G�$3%AA�nqm�*��i2����!~g"�ʴ�)���3�3�6�d�XL,�F6a�
��`@���	I �K�k7�r�1�����W�)��f�������^C
�������EiFe���^T$V�l��C̏+zj@����v?���2y�U�W�1��r�v@��ܯ1]��Z�f�;]/���4��
�%K��죢W�!@��~�iۺ���+�����g�	�%%�����m8�^/� `%�k!�IEjv��)E�,�ɱD*��B�hƢ�E��|�F~o�� ����xBk`3`���o��w�lT+�QNv�3�jAG��R��α�(�7J�"����AQ&��6�H�Km�T�G���6D�l
K�C��idQG�ry-U�Pg?�cMS>�:�R9`��vN`�وܝ�u�{99<0�Y�����$��,m�_@2��1����yt��{.�a� �ޱ���6�N���Yd����S��~�L�"�7���ډ'���K�`Z�����-Z*�#X8�&���TP��Ǉ�P��.Y�F���r�Ӧ�qͧd�����AU?� U�GP'g�{-
{a�Z;h�`dsO�Y7�gC�Z�7z�cz�����Ѷ�����K]�5Y��)Ht�И^ ?����o�e�����O!qg�+\������������[�0�Q7�4����2��'�C*5#����|�Oޡ����/�S�a[1*vh����X-B�����a\#������<f�pa�P�v���-����jώ!�syv	+�K������k) y���B�ڳ�#������{�B��%��E{L��b@��e|��_���-2F���Z�+$ �p&]-�32��a���Nη�,Ҿ�K��<��2W��zr<����1C����=�s>P�M�+q��R[�g`<|Dc���T��{��q��e�� ��x�lr8x+z�r�ʮY�Z���Uʑ�����y�@���ᨸr�_9��a��ƾ���)��G��+��k���ա�mW��`P�-VM��*rB��߲�=x��xoI�	�?�q�������pBNQ���Ąz�k��|�"Osħ7R�l"��<����;WCƆ�fY���o9�^A�I�U�zb�p}2��ʡ'���@e`@�<ɡ���Ă�"l�t8�6%��C��p�T=G�Z�����3��ůΪ�t|g/���nը:I,!=&7,�|cD�,�s� ����4v���Zw����o��f|�(|C�:\�x�)�Đ�5����*����� õ�*�`}W������з���dI?�xn���H6���>���=��3:���ķ,/�W����_g��v�����<�%v}[���̮��V>�Nv_2hc�|:���\!I(�U���s%��7Ǥus�#v�Pg��\/�ؾ���e��z�KL����>���M��2*X�ǃ��(ł�	ǋ��$��o7�\��d����vWo]t�UbU,�������ЬU?��ᇹ9���eiH/�l���=9��ZQ!<@e�Ҍ*dˊ�ќC�(K�N������3��6dʼ�&��5��י}�b	Cg�i,��=6�1"7��Q�L{��<��*���0A�l�[�2!��������'��)P���	�,}*�����\����ߦ���m'�N{VG�r����P�d��h���ݴc��������P�!�B:���,l�m�Ң�qme���L0k	�N33�{b�k8�l+��~����$T̢�@��� �]���~n��\X6�4��H(��o=m���",�����P��ܛ�c$��`��e!�|_�O�~Ӕ�$���V�1p.�*v0�R�w�ϼj���Q�1b�D�^�~:�̃1(����t#���c;3��GN1��eG��2�Q�7x�7b�E��e�l0��/I纩�����u��W���&)IR�C��t��(�� ���h�rEx;^�"P�� um������b-6Q���frI����]��0��7���3N/X����-4gx�Ba�{U�\;��#�]^P(�� [X$
*��C�Pn�xȂ^�k����b���F]x����@GƟB�����,�Ť�,�7t�Ղ��0��(_�3q��Y�Qi:���T<z� �rAb5�}�i�����rc� h5��/ap:��F#��Vn�g��H�ҝ������WK��E�+}����w�á4I�^2D��F�}�,��<N^�z��YyYh�LD�Z�%10~��g�W�Ҭ���jt��X=8��Gwm�����JZnH��R�L�3�7���K)��q��� Q=e}a)p��r$�B'�.��fß�k������B�!
��� /�^�Ae�!���׸>v!�TZ�����Q�I��.Ӭ2Pʇ�����r��Mh a��wҫ�He�scr�K%2�f����h���ߟ],AK�^�p�=D
 ��]����J�H�t�L��ܹ�䪸(
���Y � Z���nl�VH���6�+,l\Ȕ8V��ۺSQ�Z��	�q ��-���VC���8��;40y6}'�� �wid�wE���������x2����EM7A��_"_�`�Yh̉�llE����H+�M�v�Й�?���T�]�d�f3�p�����5�����g���BV?��t�]T�������{�mțC/���ԁ�9��J�����V��L�52���E!�: ��kO��)Z}K��m�0-;��v�i�;���x�b�A=�b��#��0?�������P�2��Z�"޿x�!B��fq�:3���1	���������0O�e\v\���O�I��[��tKO�T)M��=��J1����~��<���X=���,s	5�XkcJ0�Qـ���[1�	�@�����I�UuB�bb�-�7����EfP���ZU��yT�W,�+��
��sSkB�o|���Rl�!�$�	����a��M�u��4׏��5�MCZ�z�+j:��C�$����n9<ؤC)�D��)�.|�f���ZK@d��ֈ>�CQ ���5�8{�b�]Bp2�fPoF�{W�ζgYrZ��E�~���瘑ɇBIV�>(���`��Y�ۚm���QV�x?����o�Z_r\�@]��2�4�!.��~��I�_bcVr����q�5?��N�VR�F&-�O��k=�)��E�W��<u��js�2���E�7���8T��}e�l���G?>�UJ��"��w=�l�����R���M�W'�+]{:h`r(G-�Fe�*T	KE���3r�`
�d(�j�Uj�3N�<��k#`j�G�y�#&��7O�T����e� 󽃉����O.f�XS�b`�sNxWA������T^*s��(te��n�q �MB��<�b1�T
f���d�WKkC�	O�ce��{���n�̛�9�b\]a�!��g��dr\��[����V��2��N
�D�Sw)'\~��Y?�	!���E��?w���)?U����g0|͙]�����i>2Ric�@�L��:2����>�L��'�	�`�P�t �۷si���}:��;�:Gs�=UR��ܐc\�1�w%�+؁��^��F�N����N��r6	Q�WI8<&�;���n�4��|����t)YH�,Ԣ�c�=vO��Pw�~W�Vlցv:�a�m�톂19�;
a�tߡb3=�O{�Z��0�K�?�"$�Vfȼ1ǷT��?\sk_쿂�Ӂ۱.~�rM&��hN��&���혱ʵ,��n*�GX��ak
����e��M�:lJ�^א�x��ܶ��NL�2v�bֈ8��U�P���>��#��D��1�ڵ�ؔ��������k;�Z�x���IfS�8�J�^��k����M�;��#�T���|��L��;���D���sxkC�\�6��\^$)V ilI/[������'%w��l:TN�$��XH>� �x�L��'���6(�dH2vܥ��@o����VĽ� 9�ܝ)kо���P��P���]�����|(A�r�wK��^P9̎W��}�,ۊYa�-�����
^H��њ��4����p�D4~�F�F0u�;�VaP����6)T�ad�7�?�W�=�=#%��a�b+Ye��.���ί���5�P�g�͟$���_�T#��7+s�ݺ����W�8`�KZ��_w{7���,U�Uw
3�F.�|�i@D1�FRP�*,��2�8|ɸ���_2�%�?J.G�d"W�o˫	q�c�*B��\�)������$��Utk�����)�V��q��Nw�*"K�yG��i���<��
����5:�������z'����^�n)�-z��+L��&�XQoz���+���ZJ�L��&��72�����Dh����N3}�6v�j���/-xϷJS5�����ݸ�ek��� �M�`~�ʇӚ(�U�=���t����;�L�L�;��	OY�X�$ˡK��-�"<��7��"z2��o��Br5N�;�JnTъ�9K�E�l����[�Mu���p'^�޷&kS��n �,q���_nc�X|����OUwm����/�!�}Z��邔�'ؑn�L�����g ��WdqYW�l9������с_��ލ�\�����?c�QvJ�S)c��*s5ל�겅���"R]>l�ɚ��z��&�;f��T��Ax��jZ�&5�(��x���I4ŧh�U���ڏ*;�"��g�k7�|
�Z
�Cj�j�q0���=��r���������^s��{~���p������p0�7����Tܽ��k�O3��ꌘ*��t́.s�k^��q4{	`��x�r@�eG	�Fu�ӄe���~!���/����f�)D���##�A���P����!�[�� ڃ�`D��.hY'��<x�66�����N�Qk��5���+
p��y���?� ��g�g�Tq(��3r��@���8�q�Mi��z3�`�'���ƥ�ٗ�D�|�N�)���c�x3��|�- ��_.��`��	6�b)��&Y�Ր]��A���07�Je�%�<Y[\�"	MksҢ�zf�����Je2�P�ɢ��A�	+�O��C�xt<�6E�h	��Q�SwⱚI�ʙ�gG�^�t��u~Cٝ�� $�C��J?�e� ʟ[�A��	��_�c�4v�������O_5?�h?�=LC�t}䀽��̄$r��S�"[�:�$��_�r,�hu�]�u��vb�}��R�l(e/��i�2d+�/)zy���N��5r�O���P��dZ��:��1�1`���;��)w��f@[�C��m��i7�5�|�s����k��D�ƣٖ��o�k�c�w��PĴ�,"�MWT�:�&���0��wӲ��;�}�OYx���Mܠ���Z�O������#O3":z|g��B�
��C4���O�U�Ҹr�Ɏ���b5h���1P�å�U�L|U7�x�@b�^<���7ZqZ,�p��>T�q1,������GD�,��N0p��{���w�g�>���!����L��թ�u>j�=ʓ���Ɠ�`V�)���O��� ��xql5�h��)�����憎��A�Me�����59V��fkI��gs��շqM'��D{yZ������V���o$���ܣ�͵ީ�x�Y���yosW0��������}8-�C�#��6х��Х�2�Ug����"f�P��	C���Ԭ��Ո�2{R(#�z�:��I��R��jy�锪�!ǯ�{T���S��E#:�Xwnƹ"oG��n�a���S�z&�4u���)�`��E�R��h�[��#�/��Fu����
�	�:+g��A�SeT���R�S���h��<��S� �y��0�&�]��i�ڵ�?uH�����?��p�P'8H��BY�W�͂�X^5�-/D�������`j׌�@�K
�G��z��+ �����%�i�sQ,�@l�,��)5>�N���Q���oLdj ��a6��Ly��S��)C˂N]}܍K��a���ZYI�����!s����W	4h��J]�>�� �O��k�W���p���KD$V�.,�FE�:	�H�����~�kv6P3W������uʌ\�_��X�Jd��y�箐��ھ�������ʾ�v$d�:�]�1���l�z�(A��(
(aC͜�Ii�ا�����	FSg*8����;��(�L��?dX,�Zmjv��ߙ�P�As�k�9�,QՕQF1�J�A>��9g7��s�qyn.�<��?>yz�ҵ1���E�s��*��7��C���@:Ɣ�t6W��<�K�g�K	��^9h-���$��~I���"tq`�<Z��zu��Ns,DǮ}@U#_�̹�#���G��(�dF2�ӝz��7�[�V�/\���Su�F'���S��s�p�&�D2Js@�g��v���J�n^79y��BN,/joT4��{��"��]�+ƀ7�t��n��,�voٲ��|�������ؚ�L"� 7�����Bs��ʦ��(�<M�;Y�.� �g��&��;0u^��V����߫q�o�?��T�D�-�ו��8	f����V�M���3�?s+�*�]�OI�;��t��3g�0�������XO�Y�W8��_Nr���ȝG����OS�YL���ߒuw��:w��9��??��1~���ԉ�8H �V8��AO����&ĳƇ��J~������y�o%=��9En���b��آ�a���(��f�bGT���мf��L��]{nz�w"9^��Gk]U�S�ռBB��k����� W�D8S�֡&ĺ�O	g�䴛c��V�J5��B�$j&�EG�S@%��U��ބ�ƣ�EzT+�3(y�Ô<C��y�Q��2A�̊{W�X�bNi�GW����i�#fRG�i.=��؅sM���N޶�]c^&4�� s{6)~ʳB
�c��Oq�<c��v����[�.�­�aKr3�,�kd�����o�D6ps�0�m(ZZ�=R������8�@ʀ>S�"��]�A�a��]x8�
�L������4���e�B��u�pv$��i�s-/I�rF����/���_?հ���۳�ߜ����/7PrR����D �`6�Ѿ��a6����iCp�I4ƮU�P�KP������Ǉ��eN�Э`j�+u�
�(�1��+��ndd`)�V?�4�+҆�[a����Meۧ����NXX�Ȍ��aR�����e~ƹ��W���@?f���mG��	ɋN�Ҙ��@
sʐ��U��!O�G�������t���f����Vr����߯�S��Ґ�p���Nl��ىc8'O
}�ֱz ��}UD��Y�������Vr�b�n[��.���j�2�9,�IR��(;0pV��x� �+�f��m&�K�o)n���d���$�͉��­�"�j��i���]w͇���s����vT#�`:udt�o�鶏J�W����Sy�^t,�,	Ic+y�?��M]�h9Q��^1��}�&�"��v�8JC��u�?E�����w%*5w�,�991{g�.A��wh�Y�
�����.pG�@L�2^VzG`>��;�%�'�Z�I|Q��b����\�&���a(���١�b6�	�ѥ����Kz�N�4"�^��B�,�f��OH�&Z�g�D�&hi�J�7�r�n3��4��1�B}�i4`��d<������.Gz̝g��E�[~@����klI] {��5lL�\��X���Jp���T����x(~��	���� XF@��Z�������ڙ�`�O���^��+Aie�;V�Bt�C8���i?1�x,V_������w#G��x�YP2�%��|H����bX.����U,�UP*K�c�s���YS~��H6��C^�Hi�c��#H�4�{��`1,��� ���ߺ�%���v�̽��`�7*3��+��.��"av{N2�.� �a	��q�P�v��-Z��o�k+9b
c����ry���?����gG���Ú6�F5�X�߾3��_O�@Q12>:�`�p��[qѥ�8��rZ��fX8f�&�5�i!!]{֖a��� 8��L�M_r����U���-kp��o�	ZQt�$�wO�8�5V�WX��~�nT-����C�|z��ntpJ��E�0��R��H	���Y�ݔ��h?)�g`��7�vk�	�{�=!��S�� V7G�ޝ��ҹC����<$�{9V���&/��פ	֭�Y3���'H�����t@�6��T��xl���Nx�|mZ>ǎ�(�~*��Ui�0O�1���;6�k��^I�@�ځo��;F�OY"�v��۴'L�s�n�x.�L7�/����z{<~kx�%��ʹ�4+X��]��"�I�f��!>$7�'v44�[Pq:����S� �K6\`�$��
��d�0M���0̼�I�Ȕ�Y��5&��\��/y�ߵ�L����7a4h�e�9������@r0�	�k�D�Ly�A]�8������px��3gX2�.���eH-#X����x�vaV��4$o�[��U_�Z���z�Nk��Y*<�$Gd�|�	��c.�b}⎄����lŸ�Ҍt�M�?��aŴfۥ���P-�\F����p��"W�W�$ �x��|s�K�ΠN��#����U�)5��];�@\�\o�kt�Js��d��'�t6���:�l�(G%\�.al�/y�A.��
�@� �r�G���͒����t�U�g���n��LE&��%���`w���6�~�MZa����_�m1T~5S�u�udx��A����U��(.���;pp3tC�N�
�S�J�d}2u���+�*Ң��^NSj`�0E�{�03�zW�����G�Iڞ��X��#�J$q�T@Qj"��5�JO�@/~*���+s�`�'�2�(�`6\q��%�h�}�%��߄�a!ߪ��4�F5=*�ᘪP ��\'z��L�Q���}~�����6�)5TS ���I�Sɨ����"��8k5d�+w�q��؇��3?ar�5WR�
�g�x������k=3�#HĈe[�G%�h���@d�e�P
M���rW�q����i/�TM�eh��R��Z��vOzʶ2�p0���E�^���p�XW���m�I��G��:&T�\�K�R!��2a��}ێX^�=�`gZ�^Y�lD�I��O{���{m�j��eLGB.��a�xٽ0<���ٴ�c�g%�8�,u�g)�?�r��������n���2�������xQ���>�x���Z`pB�k��q�$��ڤ���@��.vV�I��?��A��d�ا�ojf�p5a �B���^h[�/U�DSKyh"cy7�u��2r���e\�Z�v��`iZ?��_�&�<�Et[�����a��?R���5�s[wnJ�0G�3!���(����*�����`�	��m°fy�3X �������m�&�^"����1ŻT�G��7� ��8z7T� �S����U9̇���n{wøcvL�d��X�r��-Rn�i
`ǡ�꾗�ĭӠ��*�̥R������z#Q��Ј�9e���r����N�a�$�� ��쩶̊���B���M�����n�SeP�V?����<�c�>�Yf���X�"�²�.��ko\*lR5?HI[9sQN�dB���.���c8���=?->��Ѷ;���b�D�+��CȔ�qm������O��֣3(G@�p�M���Q;�T'��B�T��4�V�a��Ψ���l��� ��\�
�bݝ(�j���%B��1��mS�f�G�:����<��:H�%�iBz�8�q������,���3�H*��V����A�Y��\�n��Z��)ۓ��b�`�ζ|��Ul5��t�����ԇ���D��<~���<�*�2�:��8o��%ك�}q�XZ�{[o�j����_dș����l~�M���p�^�Z?!��rp���7�d���*z*ѫ��?����EI�2�p~�
����k7��v���˾����:z���M�᳭6cl��{��@rCJZ����X:����d=��e��Q���w��.��M:`B
ުpu

'�gG�ӣ����S[�Yc
o�dmx;��a���[EH��G�H�a,� �Yfxc��,�U%�:����
e�C�d��$��&�]�,����hd���O(mX𓸟A�@T좿�B�VD��r�wȦ�	vq��,�<љ7��!1��{]h�S�z���[��4�|�+)��R-qM>�5�g~_�
���@��\0+�S�X�mL$���<^�Bg9�C�1汑s7� ��,R�ߦv��[������k*+��*f�!��Mh�y��!����A�?���hg���\��"F �<Ki �t��}��RO�O�m��{D�MlZEayc����w�����,�~�@��H��f�o{D7�a rV�n�ʚ��1�$�h��'�ȕf!����4�G�;���J-�B�6��]5�s�?ۄ-/��{��)�mZ-ǬN~�֙����v��#�M��< ��/~K�۩嶵A$;���)�y��A�������M��?�1�J�)�@�_�ຏ;�?R��\v�i<����k�ke~�	�"U��r�,#��Tణj�([�����3{�(���o�R}�_�ǎG�\.�g�3�`��f?��'���U�F���X㩕���Zﺷ�s��4��j��+����\i?�s,K�9�>���_	$��q����G������K���9J�Op�M��2>`]ힿlNhp[uUd�-���}Z����S�eJ)��M�\GjRe���s#h��wҵlh����@<����TYp�֍,���t#�v
�f��Z���1������ٓ�4x:���wݬ>	�]��͌M�$O���ѩI9[����h: A�aM,� ��^����7���f�������f���Dmy����"e���[+_�ى�_��g�x��||�l�O�,8���@N)�ȧ��c�UL��û�ވhYr�A�a�\R�s� ?[P����6ѰJ��qC/F��6N�~]V�Yo���������<+Ih�sn���>A}�G>��2�����]��V,���:R��/w~1h��s�����p���_�Nkv_WV�:�k��� ������ۛ��k�8�.?�GFI� � ��$u7$z��l��d�:�2��o LT�Z�$V��-1�gK�],]��p���\ʦdr�z?��m�,�H2�U�
��Ʊ��N�����5�Y�6k��,'S��(��J��O����Xa��-��Oy'���i`mE�%�f�&����&���s�q��t�+,�M���0`'�X軬[!.W��j�VgQ�y�J��EjK��{'�	]i������p�,J�G���n�E�2Lwl�5݃��>�⭬�{��hH�4�W�xg�$4��}@�5�@���u0������g���F��G����jh�i&�g��zG2��+����/�Z��1��]=!�J��CŴ @�(0��-��F�����=vP�`=�Ҋ�g1��g
��L�G�n���F������#��6�6(�̌��W[��K=�$�oq�N���˖��d6A���x/g���2_�uB��^M�	;�qz����N��;`�h�r��+J_��6�6V��	����
cN��e��A t�?��*�n��]��G��+X} �|���*��i��|V
�����'��^�x�1S��b��}Fe�pᥚr�����J��N�x�S)����O��}��W�B]��L\z�������[=�np��/�|�X����#�Q���.HR􀆂���E0dֿ]��!oj����o1��V��ʋu
� c�4�z���(5�?˯���w�Xas��@�E��v�1a MQ�����3��
i(|���u,�ye	�dȵ�>MҰ�:e��*3�I[���8%�������82D#���&X.J^�a5Me�����W`�Ճ������!֪yF�uf)��T_ڤ��ʘy=���\��3�b��M%�VX����rX"o��ܲC���S_'�B�'Q���f��<�lk<w6<qr��Wy��1�lH�I�k���]��p�!�ڬ0�9�_�0D��B8���M���7�|fW��Č0����7&/��1,B�Er��p�}���	A������ �O�&7����V9�7�O�>��i�r�}s9=N��͙�3�����s<����3�9Gc޵�Lpͅ���g���[�޿�oO�|2��K��yQ;t)N?G��ihJ�����Z����P��W�:M݇��#d���UEp~+v���B~`�]����GW�Wj��F��� ���P�c<s$`��bM�� B}���v)�횽\�u��T�� "'g�����w�)J�G���+�/"D��Hb���2^�Ϥ[N����тYϗ�o�ٕ��� ]G~�9]� �d���<k�RI8'XE�򈈘I"�u!��'v�g�Q8���U��|����'��Bڝ���`��l��
P��:cBag��=�����5ƀy����L�X�f����6M/��� ɇk[-�5�y��n��*�!y�}���,��)�+ғCe����u�	���n#�s8��w�%�DS���{<�?����=���QʚZ�
flC7u���2��K�OW;-�J�!Jm-J�Q0s�X�b����(>�-\%�u�Z$�S����,꿛�u�8� j1��m�8��!<�S款��a���Em;BK��%�'R���������X~wy��do%i�����e5xg�B��,�N~lȮ��t�Q�?��^��3^��%����6U�A�e���6����U\����LL�A CV�5�=�E�fM��\W}�}���Y�%c��W!=�z(G�.�p��~H��
��_b]S��6*����AyDw��`k�¡�X%�#�r�!y�� 
	||�`��&�w	VZb�����EZY������EӯJgclLXS:��l0��K�v5���.H�g�.3_F��7�&��ϊ�!�z�!Z���z��j�R���YX�UiW�EI;��tL��<�
-'%BM�a�p4�>�y	���@�"}�;���5�8Z�~�{`���T��Ph^��bÕ��C�wB���71���`�Xw�8d�S��,��%(�\xuHR]�nl0-	g�̷�O3u��p�3����N�Jܡ�-=b�=46`�A�_/qnJߗ	����u�M��Y�8�v�2_K3���ġ���9�Z��`��0n'�b#�w?���i�Mz����_-�RG���K�y�S}du�����Y���|�e)3��*E j��#8����_�y�ck?�V}��(A�ne4��:څ�&h9ɼ���6�o�v����ڗ_r:�FpZZ7�(!$�4�K��(���,d@����t���/Ű��'E"I������6P��+}A��CP�ߨ<X�)¤D�)����?�h����A�$�������yr�C��t�l�Y�l��"�j�D[<���;Q�w-��[�@��s����'�]���NN�&K�%gc̡�(���pc��ܭ�Tl:.�k���+�t�,f�;"�MF�L9ݛ�IfsG�6-p4�?�����kpThU !i~5�%쾓I���Lb��L+�i�e�c��f�훯��H\�S�O��2���i7�RX�xѴ�; `J��|�Fk�-V�-��8 ��q�9,�p�`D{�{r��wZ���vWs���enj�@���}_��ަ�+��y>�8��*�l���K�fK�rN��E$��U3�ɜ��~ ���%��w���u�P�5zaE�{�$�CA����K?O�d�4��&$E쎄�w�?�Z��Ȓ��(c�m�L����َ�ğ�*�d^:�+���&���&0=Y���F7�Z�����YL9�S���
2%������.[�Z3.F��᧖2�\xГ�=D�s7�$�֧�0JƐ�����������pf6�l�s�m�0���N�*xx�7ةe�mJ���R� o*|��Y|TKݜ{�僧�)�H(J)�{<�*o�I���w�&/��j���F�!G�?�gb}�=�S�Q�&�W�L��u��쌞�^���;V�� �Dk��S8����e(��;T����p�
�z^��œИ>9Ҙ~�^)r�wO�e�D0u����2�<��d;��N.���n-!����È��!�ś�G��~��v�I�;,� 	�{���q̑2������5�,�W��"����K���=��"x�TO����4dt��j��%���$�Æ�W2�������<�̰�Rx�&���"���0�putʔa0o?{��!�p��C�`R�²�G���P������v�7��@��;�����dAw���&30؊)c��5<a	�|�s2S	E�Z�X'�j��y.S||�Ӟx�ܫD���x�"�����f��Ix�!� Lo��ӅB�5j�H��;����%��'�����)N��R�����%�2FCe�#����qO�����?�Y�h�14�L�e���-*w]���S&}&.Ԕ���<�[F�(:�����ţ,]��yH�fJ�r�%
TQJۖZH?k9�Ե���s2V0�.V�^�>BZ��D�� �����y�����V��ܯ��Xt9֗� �x�&T�F��6��T :4���.���������J.��;W�X��=E�N$�����JO#ɓ+&02"se8����A�zpJ1�y�DPP��q'�A���m�t�_���fq�Ե�\�1I[8|Y�cۜ��E�t�H�7��&#?7n|A�n�*����=x�s.�H�W�9���zi�/{߁�	��RԳ��#���l�boQ<ޭ��N����v|,B�#�4&�{���z��4>^9զ=ӝ���9XσJE)�S�[7��
ע�T.��K5MmaGpԨ�P��G�gCR��e
��3�	w(:��� /�[��̻>�#v�?|!J��BM!+��B�O��t��!�U���A�p�¸���A0�Q�	��{f�Ͽ�/-���O��jK\X�JYU ��m)C�4|ݻ�SQ��o^��	R�'4��t�����q�l���Jt�����wǈ�9�&z��"!r*>͉����_��X� �Td�ɱO�K�95�&��G-���R �ܱ�)�gEs�Mھ���3+�6^h^��$���H��8&��S��4����Rp[{^Y:��b�~.���)w�eݵ����TR��R 0(S�ʍ�'@��lF�y�^��� �We�;oւD�f=E��ݱ�p�Ѹp/,��+�UI��lR����K����t��굪�3���,�������;�zX�hp��˧§��J�+���0�b�X%���X����6���1���A���jC�*��*���n�������S-q���
�%5�t��}�4WU����2t���~�F�K���>ǹ��x�&��6OB��廗%c?Ȱ]^�a��$�^k����H�y��uDG��q�(.�i4���[Z'�n�U�f�rJC͓���
X��T�u�'4��F�@��Z��*���(׌���wq����*��㢝/���v���Hπ�½��$��tV,/K��"�[�1_h����qlZ�1����8�i�*���bl��Uͭ;j��ag'E総�x�f�hǒ�2��	��G��&��,Ap�M�����������k;�����n�j���bS��%(,�� }6i�0+Pjf�l��nME��!��r?����,q��P�w���ί�M�ӯ*����^)�$/���J꣥�i%K�fC��Q�J���X��5�כ�u�{I.��т��g���E�v
�DF��i�
5�`$nI��7
��ξH4-�א�9-a}�^��*%~����7)��7Z��1J�E�4���WB@�����.��.۠�|���D\�lVQd`����(
��+�7��ݐҕ�4�\jH���y m:UaJ�]�_#t^�*�yА�Jo���S{+�HH@)�ޔ�l�R��uHFE>q^+�v��S���������1���V5��V��x�C��0���ٷ�	� H�cMぁH�<��>�g�1�hE|,s��Q�J�ϓժ�� 3E��L�����r�w����bS��&P����O`*���L�<�|�Br>�E }����c��E�I�yB7qf΍RE�;�Cj��nxs��/�ؼ�ᚕw���s�"��H5s��
C^^U
�8���'��Y�t#� {d���E�;���`�?�u���0����pM�r�`����S��3����?bۮ>�M�*���\m��8˯օ��)K�3�?�n	������=�y�y%���Q������$�a*���&��)��?]�U�P�0v�w������&���Ĥ׫���k%o�����E�-(Qk����"-,ohʚ׭1�7��-���9�ֱ]6�+��� ��}c�p��쑉3�@Y<���/�k����y����9�i����V�*�삙a�P��#d��&5��qB�3llu�D�����Tg�b�r�,�$�Gaa�N�"�gw���V`hW<����|�&sR�ʄ��z�S����A��?&9���p��c"���
���?ďZlM��vV-�������2#�9_�ÙM�U�P��6f٪=�χ ��f�f���8o8\d�_�Ǫ�E�֪ޖ6��c%����4�v�,��G����L�.2/`:њ�+�;�#�{�_5�m?9���ax(�����8�;)����?�~U�U]k��=�\�# -N6gc�A��a�J��#h�߄g
�[0��[Fz��㋁�2�1Y98V��R{7���W���9�y��CZ�VWo�t|��d�VK��Ya��/��}��([٘�EƠ4ڴ=��L�j��|����:�/:���'���<m��k8Xr�H��{�=�����:��Y�pW `�v:�O�؋TxW���Rb�n$��>�d�t+�(�z�3E~��7�t+��}��{�(�w�����;UP���B���я��ȡF��#�x|�/��}�2m^����_d��'�+��Q �Nf��dOb�����$D��
Gމ�����e6ZY��i��Ra�"�i_��!p�م!�j��2@ݤ�
�)G�FT*�[ԍ�p�U��Z�V������@C)�'`�t�Ir,����}�Dd"��PM�Û�e��.f��G?�Zn���%9�I��'�W�P��!�.���\��w�J�k�h�lK��dvJ�C��'�l�lu� �
;F���~'݂&��A�eoIp]��9&cB���J��fc�>�p���R� ���;3�|
��8��i���ؼ/������ӊ�/�;Q��+�U�1�[.caqxN��P��o��c�G���e��Aw� �{u��7�}+��Z�U�	��� ��M�5.� ,ǫ�#���oꮛu�{ Pc��Np=��s'GL{��F^�(D�AV}ǴO�ȷ��@J�݂�W�KF������kb%�����3��J�)�OE��X8���P��J!=�W�����k���ж�GS-�ֈ%{�,_/�P���:�p��f2�𯝑��)/rګP}�KweD.�sڮ�3�X�#��wL�ݚZyU�������_-}@G5��{��hV���ID�ӌ�q�X��qs�ɱ�[���>��Rt�~�K���>��x7�ˢ��Zg&]]�^�-L��o;܏�=��E�H�^�I�Q����y,�o�,V��p{jH=!�儓�r�Cav��?�s7,�u
jX�remD��}Nr��h�o�T;�~��1�|bc������	��ӧ�p��~
��/�V9jyȃ~��Kґ,�C�ט+���ew)� �|�r�d���+������dA)�S"]@����7�s��OĔ��P'����O�mcEX�C�o��2�mC�MÐ�+r(r1�I4���^\����������3�<._��U�9.�Y���}!K~�Q��밼�1Z���c��S<�9�̹&��6��ϐ	��)YE=���|Ͽ�o�?]�·���)�p�������5������2Z��a8�T	���:s�f�}i�H}��6�����)��ʯ�V�`�%�DH�W���S����,+83V��8�Te7����ǰ=�#N�&γh@��c��ޙ\y�H_#D1��S��GGĪ��1�޳��JZ���go�WM�Fv�A��E���_�����U޽V��cbG�B�к	\ �-��~�20 �m۱���,�I�c�qi����k��
���o�+�\��*���k��Z�� ommC����Ӫ�����ƀ
M�G�Yp_�2�Jt0��cĵUU�}0I�PQ9QZ%����`�� އY�?�?.L�9'�F�_�$f����6���*hae܈�:|�J=c?ˊ
���xD{ФO{��9��{b�#�.�n��=P��|�U�1�1�ƞ���a�>��%q���p@z��}*F���	��siJ��Aܫ�Quv�����Cf�+���ކf7:j���e8�5� �Em�Y<�Rt�O��\�7W����z6��h���0��GM�'a�z�z_���ZWDK-�ު�U��ЬZ��{@OYĒW|���݃�D�)Sq^��f�$ɻ���k�k�	U:S�ĭC�-�#�췳��\�l�{b�ns���*.#���� _`�q�!����L�G,�r������@΋^��~�\w�����		8�Yw���@ޤ�#�&�|FPX�,������n/��/j	m��
�k�k�gX�/4���D��=i:�q+��� �'�BW!<�!�I��pG�<lͪ)Y򌍣���L���я]���ʔhR��'���k���ʚ���9�L.9@)�A3��V�|��*!vƔP�i��i��ǥ��b����="�Dd� �ۥy�
��q�a��>��g�vH���WΗ����g��� /�ל6� RЙHN��M��v�^��ЬK����T���\ث#ai���7���Ҋ9�W����ąVa��xR�Ԟ�~�n>p�f�DSpM���	���=���v���f�{m��d�c���x�e�6�,�{��-f;�)�?B�.�g�%B�M��9 �d�.��h�	�P����l[[�)e�[�*�𹿬��9�۪<�|N�;�"�'ܲ$k�,�e<e�A'0˽��B�?��a?�*�psg�)z�p݌R{�'_�62y2*���#D��A:u}T_]���$�P�#����w�V�� W$�qg��o�^	��|��v�ϭ^#'�Ч�yo_��z���[���>�h{�{�[&R�%H��
��	��R�yA�T��%~E܃穳�/8�baC����9%9�b�"�{�n�/oy1���GmY@�j5���VMa���F���S��\����UbC�wM���:e�M�C�$!F��>��h��i��:u����헴۽��E�_��k�?Flw*u��V]���"|�h�[�O��'N��e#F7q��C�'��m���({c�x:�Z�c�TI�e�G�8�a�{Lg�D�Ƥx7��_�B?���9e��n�� ?3c���@C�W "	��ŒV�d���u��PU��\Yt�'�-`��˗Ї$w���*aiI؜��]>��D�Ͽ����ɿ��u��=�P#������Ð���M��W0���V���ISL�z:τ��.R�>�K"�O�k��&����M��9��T�K9�^=�����A���>e\��)�m�cu9��>��oY��n�S�f���P�3:����-
N��##Բ]�\t�2'�Х�螯6|6Z���?�[��<l-i�ls=��#��`��9JFw#:���C�C嗹3�������� �i��:C��{X�L�h��Ĩ��+`
P�H��)���H�~�|����CG{�v܊s�y��SD��7	lX����>��
Y~IU����{a��*�I�,f}O�$Zg�<K�!e�� ���ǥy��}No���(s�k��pr���9o
%zz���Ƌu�QCB���
�C�,�(����m^��2]`Y�q��6�,Z�/�������(}b�%i�b�){5(��/De%��A�����5i���$xK^�~���^g�h{\HY>�.�ˀ�
o��gN��a������S�ίK����݀:��s۩�K	}q�9�M��D0Y��tqi����9i�K�S�ʛ�����!%��p�bd�2J��q�CT�v��&#�P���*dq͑)9M�v>X���K����V��'�wN|6�#����Qڒ��o1T���gk-�?�3��Q�\ ޵�
�ɖ�8�z*�m5��sWeހ�$����8ۙ�}j��;n��������M�.n��[tc�+E��$@|�O��?����aEw�)h.5߬��¡6 �U
���t�j���R�@����<0��,T{u\`2p��I4/o�-���tG�
�7;���E[	��2�#�~G���F~_Q��LJ��}ZY[?E')�ğ��^��?Z�v������_�[F�,�kXM��4�yx/�M9�#zi䳴�����"Wsh1Y;�2i��WE�z4P�;"r�i�5���0�:��|`�T�X�T�7$}��"�-�4�HV�K>�X}���Φ�$�-ػD|���gk�ɓ�{��H�y�����������/�3�`��r�F�b�[~����-����z�O4��B �b�m��������1Z���ҿ)�In�lA�?!�DO�(;~`�$F&�!���f���@P�.���^�_C���N�޼?@�~�"��"�5��<���Um���&�2	����V�k���<ɨ[?�h������VY?�1G%�G�h����z��H'"�T�p��K�i���1�Oq�ƀ;���ao-�s�NO�c��BS�p�ƿp0{����S����x���a���,y�ސ �8,�������ډ��5�G�}ܕR6�8����I�����K���U����bڙ;�y6�O�mWfgmlhh��]O9r)�Do���;��?�o���{T>B�#��݋��qNT�ĊS��Ycx�P�(�I-�8��R�x-��UmF���w���׹��~��F<���p{��9~6~�oI�����L�^�G�����߃{dQ {������=�{�39��k��>bgq��zz-GU ��ش�\���J,��5����\�\q˔7��w�i�/P�^��)��'>�1;6xz�+/���m��אHU�^��	�ӫNS���5@d�"�$а�2��Vha6�`f�
�S;�wӜ�`lH��p�����P���t��T���i��(x���3�,_�r����� ����OG�ݖ���Dk�8+����XĿ�H�,�����˥��=�q2̸`N��yp|��ߑ�/xK�yT���`t���ɎQwک"��=UT�Ө@�� �W�X͏5��L.Vu�j
�k�Ƈ<����iL�eв�t*�с-�?��)���Q�a�j�K*x��6���RU�x�i��=+�V��H��$��<6�gb<���"x�=?�����󮒶���qΡ�*�7)���`$���謢:)gb6��V�ZQ�I̔�0�O����j�o���F2bL�OmD>eK!)��I��?�#��I;(]4��%<��H �^P�)UDT��V,���ֲ̉���7�A�?�w3F�: ��m�� ����%�>OP�EB5t��-|R��H!��z�b�>U�D�.��=
M�l��z%7�;fѠ��ɥ��R��-?�M��ѽ�>�IMg���l7��	H���w�Î\���gS���P��5���@������	�Ѣ�� :��<D�f��۱�UotKqL�JI�z��鐊�+�� ��5ju"���CV�9�Ȃ�����j(XH���� �*c1#v�L�_���i��ݣi��
6��V輻*�`E1m�3Ȱ	��y�4>���X"bld�[&�1~��ts\�>1$ �%���D�r�t��˳���Ł�.�]f�ˎn��c+�r��(�$l`�AG�� J��L����X��t�ͻ{ m��g�&��b�����3�"pziͰF2�n�AjCn�O��Q��s��f���c�n��@�x1�1u��YjOd��������7�U`v��~矺�Ii�5�M�8{4�OڝQ��ڿU��l8�gv&=)En:�>ř�r-r��2iG�=�_Ha�!�G��bL��)#����+̍����b��H���o#爩۪9;�߅I6�?�@K�O��Ĩ��b9,��u�߫�P]�2oY�M[&�xZ�.�a�ۼo3��yt��}аG5D!�ȅ=�3��a)P�;�|�u|���	�6�6�LY�g[}���rJ���K~q^#�k�^#�÷�l4�\D��X�ʒ��^W���Ʈ4ې������b�Ԡ9���v���k���d;��kp߫V�M�y�K$��=$���uj�3��|q&FZN
����2��ʒf!��?�"c��L��J]aU��-���M?Z�O�5B��D��q�W����o��* �3���WԻ<������𠫆���~S6*n��W�pe����(֩�Coæv
9���N?�h\�N�;��e��T��§7�<{�z���r�22�6�{�[Q�8y`�+�s����.��n������ܟ�ߧer��uF�?�]
KPRoO�!$ú �+<\۲)Y�5V�����ľ���v�:p����ġ�H�N�j3�­����l뿀V�k� ^���_�ⴗ�R�{MQ���)�-׵f5��.ي������n��#�ϫ�q��}��MT�����]KH���h����8�$�<g�m+��߈�E9
=黚�h��|�ɷ˿��]E�o需*�g0o�9JzJ�Zj\_��\_�������8�\H�ѹ��g<D�c�0Rw�"�Xhwc�~�ێ�+�`�UQR�hƾ�����qy�Ļ���Jע1ؕ�'�a���'���2X�QZ6�����G{���'�
��3�<�1��o"[��E�md`�����O9!�q���'�C!^��Э��Ie���zKH m�9�CtUi�"2�@'��c�����I��΅j<# �3���IW���Ն�mD5���j�f��zz��5�j�-Nu��R�+������q��$�)�oCS��tY��y2�Κ"�o8|���0(sA�7�"[�J6]H�vu�%s�ly|W,gA����5��-��P��&L�z}~j����UQ���o3�k����&��GY�x��y���i@v�z8�Sk��Ds��'H�aYh�����Nٮ��F�C�/�/|!c���+#��E׵��,f�' �R�������4����ԕ+�:����ɰ��փ�+�,|0@���l]�Z]�Y�{�[����ta7t�a�fZ�!�����h����@Ae�� �`�/j��8]�3ٯ۩��{2X?��4�����2��գ�ao'� �g�^��@�3��p�"^]�EQ���u�:}˼��5G�^���f��)��a��n)�}/w�2��aÆgVP�������j�J�/��t��?���|�P��ڔ~0���@�U���`�I?ZfF�1Tv���`�QK����p(��1y��s����pq�P�h�T���$���a��h�����%�J��B|�uq7~�Հn`J�����S��[��f�WP���Z�Rϛi9]���� �w��®
���ɵ�`{�B������~nEj�^�?��s3��	�W>u�I��Ӡ�/�|��\ �����(���|H@��j	ό��	ޡ��H���<T�|�AV}X҂����*��;h߷���J���?���a4zE�-[�>q�{5'X6���_$���2hL'�2OVFK���{�/�͐���"⍐��ھ�r<���* Ŏ����-w�Y�bJ}v�u�%����0���;��7Ñ�V��74����+�9)KARx�(BWk�m2��g�E�!~��r\�mGw>�/����UH���u-��q٣��v�?݂��(ݱ��t�����~��/A�͗̍Py��	�[7� �ֻ�˗D*�@[��Ó�h��wf�{��@��vc�S�k���l����!���Ė��R+ �WQ��l��)�*_�<�n(��a5�A- U�q��5����(�&�iG�Z�D�<��Q���
J�F4�nP���i�J�f�j�Vs㑛e�9W4����j��?j�Ӿ1�(��C�oɀ/�TfH�]�݀�<#y�;�	��%2��ޯHR����(`iF�R^��n�V5U;�b��J��#�"�E42��3#xQmHH�E�K��~�Rg�S��Yw�d�Z�����	 �����@J�!���iS�F��b�5���(K�X,ά��`���g�*�ĵ�3+`x2��� u�'��M��"�Q��j������(�p^Â��5�2#���^Y^���K�c�0��'�\#�է�t�pQ$1�g��ۏ�h�ل��َQ�;��A���ń�wՁ�$�	�h0�t���]pP�I.��������h}���$�I)�+�{n#��Ǳ�а�aX
�`�O���5���_�lgԿ�����)����^���Ni��i_b&���W�7�)�/���
��~*�K�G*�Ap�¢,y8����##��х��Ud����c���plh��P����w�^�;���v����kH�uP��L�����7�-����%��4���^7��	��w�JB�g��:c�#�dm �BDx��f�!3���aB)�{=0��&YY�c`AbOq�'��L�-�v%�O����W���#� �G�\�v�����(\;��g	V�,��#��\m��V�E]�q��5�q�5/ʳ"b�5�t�7>���߹�f(�y��?��Hx�	½�F���q�eo'X% �+����l�u���Wi��L� �&i���֪"��"��'=����Z�"�H��7���O��#:�B���)
#��'���2�5�G��D�K�x�i�O力
�GdM�i�?��t��ة��j�Cay��� �>�iak1��ݓ�ĕȝ�	����<:�<v��>W�D;}��w��F J<�G�U8��3����B //����v+� �"죭Ü9��i&��� ����v�n��p�6�]���&��oE
�*!:Z� -�ԓR�5�s��w�=��XR�n��dc�=��9<��b������?yz���9ʽ�-�%�,[�Hl��U��S����!����pMn
�!�'Y�!�8����͍�U��nA&bئ��g��a����0q#`;�����^�n�@�E��65�Ͽ�B���ºvR���8����ש-���݂p�2�G�I�}��vj�R"'����{[#""�.�s�H"=m��U�*<l��6ae���6m����e��!�
G 	���{���y���|Y�k\$�-'a�O�-��踚'�&t���̑�J�?	#�d�D1��HUp�	�!RCO#	���3��_k	�OzJ��<KtR�DQY����|XQ����u�� ���d����d�y![��
VQB ��p׌����k�m�/�ѣe��1�-�Y7ďF҇gg�-��"F�p��l*:�fO��X ��!n�EC	��ٞu����ƺ"�_�B�O�JKy`��;=��\�$jU!��({�R���6��й��&���RwB�����0�r�w���$�:�k��N���ml9�i0ab7�b�5���y��/jl��7��f�ߟY�rbFN�j0�u5�7nO��ZR�M�z�F�u�ۀo�������:��t	�2�\��d`�<�5��C:wL�?I��q���u!�;���~�54;��$������w,�:�ﯛ�6q6I�9[	��ڒ@ҋ�\���PRnE�5���Y7�����ڏ�m>�/Y&�d��l��՞p������tL��dL%�R���q�Rc]7��hB�ҸK\��|P�av�?wt�t�  �����ЦݿL���h�(�o���Tz�6�S����Fc�K�,I�5�7�.12״�j7˦�)T�#�E�R�!x�x�N��SV�n{-�0v�)�%�r!b��������r�������������q�s¡�<�J^F�S�l������]@ma�v�W��1���}崵!�n~M��֢��{�.���Lѣ�/m-�W�P=�s�ۂ�c`���3��0������)���/��9�)���k��9�CQ����m�����!p�(���V�tM�lh�G���ND��h�*u��0
����0J,�B.ˮ�Q$�%u~I	$��d����,nhi�7�����B}�y��W���]��]� �k*�����@��!�&�pQ�^��G�<�o��x�¬&� ǰ7m?-����D�N0g��y)#��҅-�7E�����ߐJ��F~����zQ���KTj��H݃�&T&�:��m:[V�9����(g�E"��ȵ�V\�-������u2ӗ�����ts�v���e�*�A\�*S[@��69j��3�H����7�UB�3Y��	
��
��ԧ=�F=�[Q�̢׆]3�T0CW��lĳ��ɓ�K���&>�8���aj�	�#v:�N���i*�QJ�����݊\����GvoZ�mv���p?�6DHGrn�Ztd�M$�?�C�'�K�A��̔`�Xi�(�B�fd�E$�.!��������;H�96�*�ʏ�ZZ�i�|�Ï0�\�:ׁ�볯2�7���K��WLua�@��Һ��hU�����~l��]P�������%�3Qqd�{���D�X<�Kp�/����0c��0��vB�=a��Y�5�|O��P��� ���U�!�nOۄ�a�񭐹+yi+���}�i����Y�qp��|?���NNR�WQ��e���  ,�Bʈ��g�Ɔ�FZk0��K8~|�#2�n�`<l��+�'u�B��lN����<%�<ބ$�M\I�@l���U%�e�B׌F#�Y�q��{�'.���;���!L`��D&/ѝ���űr��@S�e���WSԭ���P��@VA̓n3�vAUe:`��6¢�r���)6d4,�z�S}#�hK�
�D�"!�8ȟO�	��mUH�"���$û$�m��xB��<l:hD�z1�4��4�̈�0��F)�"K��gS(���������\��Ti��hȾ�Ġ"K�W�^�t�iJ֡co�
r�˭�K����'��Bв֦
�x�k�/��
7R�Ca=qC!z?'�tz�v�'TP_b�����9�����2��[���ε8��d�H�x���u!��W���O����;4o��k~iF��i��8��	����.^�^/M���:R�O�
�?	u�YO�K�*���C�;lV�eq*�}ŧ죸�;�-�sˌ��Kc�Z�uU�,�߃���t�i0��7�7N7�8Wk�6حr*Q9[�Vd,��<��~my]��ۛ>�*�3���m�I�^����� 3q�:W��&m,��xg��렛��a\+�G����㔝�h�#��.��J�� ����T�N�;�V}�U׹�	��=>Z2�1����u'���^�N�U��<�t
���2VƓ	v�n��r��E����u���֭ZК�oa��C�n�&�ﮚ�sBխ[�J�ʥ�
.W�����|�&��f�_�c���S�p+xE���@o��ב���=i��A*��wS:�Onw��W�B�C[7�	���ܻ��?���#�K 9�odN�m��4�6���� -g�g�h��i��(*�{�5�����dD )�%Ȍg"����l�����YM��<��:���ni"
�qW(��_�x�${�k?σ�2(�6�&妎�h�v�i5�Ay�<s�q���&@���d��?6��*���!���ڷ�j�t���s�`��2�י\�s弫�W>PV�/
EqО�������CX �ȗ�Q�@�-����\?W�!��<n�6����Г3�je�ē�`���>o�&����7��IJa,��X�Aԙ�oL���x�?݁���(:����Lv�����Q�����7�Z�S�`��g4��wq-:�E����8Y!=U�z�k�2���ȅD�	���<�A+����z�n��V��]��[��T��EX$⣺�
k��L��L���9P-<e|�M�����W�?�Ǡ�|��k�L����|<�W�
<IK�i
;(�0���`����<ֈ����^�����9{�U6R ጃ�̦��b+_2�5L^��=x�=�V�ܕ	%ƪKÃ���-��L����دm�/.��h�T��%���4_���U''A{�ڏ�ǝg���Z���n���w��ϯ�}	��y%��c��G8�t8-�K�&�f�l�<^�w1��M9�Vx׿ǽ|<I��hb�M�C ���?u�Wܚ�Iry��6rh��fŶ�{�Bb����%�QB�5_u'ln?�D#��xYg���z,�� �j<%�AE ��TTo��|��߲�8�x7Q	)�K�;WT�AYݘX�9|����I<�Vjg7��zo��p����M��ҳ�J�����uS��3��?�.�6�ċa'�s��~�K�de�&)��k�1 ��/�r��&�Ef$�w��5�k�����q�4H��:J8�y����~7b�Z�_��:OfF���(�Tz/�-�>]�=��$cx�_5~�P��ux7�Etr_P���Ŋ������.�U�|�S�Lw����?;��t��dy���G�w�5���`���#Bv�����Rs�a˧u��GCY��r�p��M�n 6�kO�{�dt{#����0�g�Z�-��p�7}��b��-|��AYN��q�Ol�(˄����»d���M�*��� �ם�b�R��uo!0uθGb����������
�S�٬L������v����ѐy�kW�Ko./qV��× �pve`����iK�J��@pU�@s��;_��pr+��&əQ�D*�I{����s�e7��=�;s���m�1`�O��� II�X���=�����9鮵��B��sɫzJ3�𓄷*[��d\7�	���O��8����<�-F��|�(�Zo�m"wO/Q�����%WV��/���&����`�\~��KHǫ]�I�)�s� fc�'ഞ�A��=�&;���~J�2��!*Wo�T���	d�
ޔ���W��y2��W��Ɨ;�_5_$��Y�:�&�RB��D�}{�M��d��L�}�@���3�"��V4v�Hk��u�L��zcd�ʜ��*��w�&T�	���C�˰����w.�0(��GP`%�퀱�"�5������ �*,FNS��W�7���}"�~RƇ׼��z�k>��3��i9 �fm����/o$�oE��o�#3\�K��;�~Ȟ�_�^&�I�H
۰|Ο��z��G��A۴�J���4�QҊ뮠5qvsB�k��E����z�(Aٲ+-3L�PM U)�ň�>~�J\A��h�g=�-���v^7������<�-a�C۔_����*z:-�j��RԽ3.����Q�ھd�y����a��:��0�=2"�� 0�^��V�WWj��'Z��`qh�Qh2?$�`���W
Ng��b��Q��Ҏ���0�.J������H������ty(Bel����:�KQ�Q��+1�T��8����\�����PD�{�X%���[vm����J�>��I=��x^�E�s���k빓9��1�a�#Sx�z���L�� dtd�!�ٜ�C��g�n�u� _�PWE��f:>A���ި�]"�yb�� }{Z���\O:N-wWdT�N����pu׺�j�?cǦ��Ȕ��-֫��;L��Ay+��V�����%��zL�����ؐ�(�����>�;C=�><�xۮZ�w�L`�����KA�.id�e��O�?��%��=��?Hg����N��w�Gt$���?��x�2ƾ�\⌗�HmU$=��/�����d~�	�	A�VA�L�p�p�C�������*����Y��	��?b��Z�+v�����hݝ���R�����j|�e��ZIF6A����?ˢm����E�2���da��u����pMGkf?U����U��UQ��] P��cX	�عج�c��4V}M2��j07S��LS�@;��-Z�ٗ���r�^�>�/~�	t�S���\n��1�)&��TX����o;E��_��s5O|[H��՟����>bb�9�a�]�Ի󼑥�$�;��ā~�L�*�B�%,��B�ɽt��qx�J1.?���+ݔ�|�\p����9���"�:/E�̴?J^�)��N���wg��:QW�Ī�Dy��n0��6���n���Y�@1��:��iس&�P�wK��wW��Ú}�$�{��(ָ�����bZ5�L��B��q�l��?��-C2��Xu�L���j���|����2�Z��͎���S~��C�7��ϊ~_�z,���C�;��ntaG��E$�����
(�y
�H�#��4�Zb#W+�[�ƻq�ď�����(��
�4S��(���+�ߺ�%��-g-��,ai�h��z�i�A���h4걓�s���r�Zw��St�mJJx�oC��T!aPo��[�����k��"�  d��Y�󭦤��3���Ri�nF�6Ĉ����&�:���k=P��I���Wo����ʸ�>t::`�h^Ρ𥢧ܶ��p�| �v���Ə�r�IQÍG[8U[ݭ�:�r��N�g��ﯲ8()!�����YF�,(�Oϐ�3����()GV�K�߅oT�3�_r����CC�|��*<�E{�3jm���bg�[@�l�w&��$�2� �Oˊ��" ����5���y�B���yWB�,S&~��G�A�'�l?�h<!��紹�SA��TP���q�)S.�ngt��	�:kv�/L�1j��O��/��I��7��I����Z>�N��)b5ҧxMn���sj�?��OY�l��&S=����8��� |�!fa�?������$�zM�|�O�{�bcu����˕�Y$e}غW���Z�П��(�R��p��"T+i���V��oq��IŶ|��Gi���i�|6�?��:{>C'�*��iL]Sg��A�7�O����2od�=4�q�|ۗ�?t�q��?���k�$S�8P�+x�%A}gQ��� ���$m�������z�\SjL�=B�L_S*������BH��K��Yt���x�n&L�7~|�dG�T��wb�)��5}�0^'Oh���am�U�-�����8?����G�5���y��k
���j{��2����~5`�H���d#Mx�6MM�=M�5������q�@H$��-7�t����T�ˢ��8��� � �OS���ꎉ�t�ʇΫ��3��yw�_��j�?��eѡ��r�g?f S�t��j+�i�K/�"r�rj�������wc�x	�ݘnXi'Ά)-9��8
�9�g�/a��ĴWg�=l�rM���i�[���q�fjy�20����l����ݹ.q�q}�A�癣yŽzb��~ja`ql92�	+C�gq�k�� �m��I�#"ô��3~��Y�Ł���k�p|���Ჲt7?E>=69�in�SU��^3�*F��ʹݥ�#���)9�B8�nZGf�ɤ� � ��w��amy9s�3o�]���T����-�]�̮f,�T(ǚ^Tg����S:�9$�~ �>�M��|�V��o獫���@�f�G�BRfa���NH���΀$ ����`��@��7�%��#-�΄ *�n�� ,�Ay�cSWl`�t�����("f�pR� �����=��({�T{_=&��"V���d*0�����x�����~��P���:�%�)g�?7$CD3,��%Q�K5yS��`���@'�Y�d x�+��]êqY8)����̫���?�12��|�p^k_}�]�N��ʷ��
aD3F��V���9A�JYִ)K�����~��E�k�#�_j&�#�U��<�ތP�/�@�����B����mUv�sP���ﶊm���>�QT�tnN`�SF ��Pm��
���If5�@	����+�r�tў5��T��z$��������M���|b�w�tA��in>�z_�H3s	��㤌����0���L�@�f�(r榜�
�(C��Բa
�yr.Z�iё���_q��e���0�����,߶�#�a�_}l�&@ ��C���%��E�/Y����&����e���f�=�KG��t�r��19Rg*>W+�⛺����Io�&�mxىy������-孤�Az{��\߀n�_�8YI���r[vU�H���~}v�+R��M�|��	H�ׄ���֑q�J	}��gv�aXq!Ɣ��c�=\�Oٛ��o�o�(_w� b�E�����!"%�*xf0�G��d�ɀ(tRU��ݫ����RM����`CV��v�B��O��O���� 5��p^�J9�p�d>*�&����E�����G�q+g��[�%eb�y%�0��'���h=��
��� ��\��7	3zQ,b��"�DBp1t�_/���!����F�q���"!~�$��ZN�Fƪ@䕿\�γ�����Fn01��E�)p�Vq2�vx���u�>�	��fc��D>��ݓ��jO�)_���R�`��H��: 
gY����#�J�킢��3� ����$h�ߠ����M���$N��N�LǫIkb�^�2�O5�������t��U�F�����z��·6'w���r�B�^)IJ}��9�{/���k	�.��`k�;.�zK���Y�Y��F��B�`[6tH@�A�ˬ��F�"*ͪ�Ϥ3'w~�j�����\$���-V��� �j��.�k^s�;޸�P �M���K�+�_�ih��Vq��=Bw�s��X��Q����D2���T�7[�6l�c�Ia��0<�Դ� =������ɧ����u�)��t�	]�r�-����c�CKI�%��n'����0ܢ7yo�8]䞳��g?>4�k�M�=�l�g� ��,h_���	mH�cڟ�����:����Tdh�d���z�rE�.��\DŻ>�e ����	gl�ƨ��.{d�`E6%��t��G�H��,�;Q`�K��e�+b�~��R��<��H&�C��N�{ķ�z}��˓�`߬�5���N��Fk��Q�/�p�Qjb�S�f�R��O1t�u��S�G~�=N`║fw��9�R$/X=�+Ʃ!�gq5�A���-��h��w�G�Ch�{+��
�a�y�Z��@�e	����5�	����]G���킚/�H��ۡn�����b��.���<42U*k�,��X��n�Ʃs�ᵛF��6�z�f+R��O�����=��#��]�D>�2Ǹ�b�AN�ݐ]�%)�tA��9��!�b�}:����OX�9y!e�|�F�/�������I�����9O>�
(�5���,ڋ<=er�`�T�b���P��G=�ToY;���U������M���I,7���urd6�>;�`���#�~K�j�!�'�j)vnR۱7`UmҚ=ex�/��s�����<�њ��Ε!��4f�3B<���)���_�V���^<��������}8i�kK�Y�$��}�%����`c��3�Y��y��L�4�<�>�e��Wq�E�=w���R�l�	b,�\{VtN�9���&�Oc�3#�xz۩��/��Owx��_�'��|���2K��W�t�e^�3�Mq�\�@%��4�&3�f�ܰ�Y�b(�g&nn�8N�.B��pK��cl"�d� �tB�*��u|��	�i&�h�#���>f̒W�u;ա���W[�ʵq�£}s���>�\��z��1v	L_w2����J��Lq�j�sF�G��Є�G���Uu�8Jo���O��׶��d�^�K|����1��ci>$��Vw�O�|��|�����#u��8*8f���ԋO6ď޺�Ph���1Y����7��V�2r�m���;��Y��4��4��4���@eG��x�z���L~�` ��+u3Oþ�/Vi�x5�<&���O	7m��.�-x}�7���A� ،0��$}AG����ǙS�юNͪ�J9?c��p?�*��]��?�L�P�d�5�v��M�fF`��O0lW2��c��k�M�"�[r���F�\b����ބ��|0�T+QkjtgH����k�Xb ����m�h�T\�T��m�v$��R�U�+3+ي��8�:충�rY�U��:�_�e��/f��K9_I��{�Cx��9�Q,��[@���k@DQ�%�:��"wC���o_fxK�Û5vD���<-��12�[۵�r蓞�6�H{�A$�6�K�O/]�o�t�-5J7C���QOc��nb�bSQ�Be���A�zјKs�>/&��iU�ڴ�ik<d����U�-}R��Lb�$T K��cm�uզ�X���x�gu��⬸��1j;����@�c��&:���Y�����Ac
��$�S�U��=�r~�i�ǜ1e\�]��Z����3�+"�Ke�t�hg?����$T�����?�C~��F�W�?��Dٲ"���{,k=]lKj���)�:ֱ=qZ6L�MzV-O���cp���~�0,��֭~v�/�w���$�g�D��7�$E7��}��E�V'�P�18 �rx�W�=��#�.�MFX�H���!�"ӣ��b@L���4���6n�8�h�n��
x(<�}^��h�f}
�z�jy§����NW�(���@���_ց��p��V�{�����⏂��(C�u�X��p��dn+Pn:�����+c�g��씞x�Y������D�{`2��J�����b����'�;lr�M5>ڈ��ݢ��=?^��?-���k7���`�������d�i���� ou~�����-p4���[p�1���
�8�[�� +s�0�P��ƌG�1��>�\!��f���B��ʓc��ELyJ��8❫��9#�B^�Y�O�6!od����_PF���NM��P���%�N�_@�Նk�����Z�S{�@6��-�9�E���U~�>H8�G\�Bg�_~��ط^��� ���atB�w�U�/���*��*�٪��D�n�]�e��?���\QK�m8E�`&z�ݪ���qWɅ�vz�����Ҡ6�K�2m^ogLљY���
$>;1�_d�*��w�s��&��O�����[&��> 1:_�E9X�v���Z�̴.0
Ɣ�������+�&�ߠ��`�2z��.u����r� �G�t��sG�ss���7�c��X��s�_t��/�J����χ.�&e� �\ئu�yh���]�F�Ȋ�F22>�<�]�5�)]D��͢=�� ���D���W.�v+'J5w/%��!��iw�c=��C��Hƹ�	�	�u��@��-G�>N��L8��3u�y�tn4�r��]"0�W���GU�B-��"��r0�IU�&�;�^�wJ\�f,l�Ǿs-��Q ���9�>C�E	2+�����Nzy�*��J,�����ځW�5��tW�.v��a䨀#>�Lm'�5�\�j�>���W-��ֲ��v�ov#�?6����:�8����{X��Gr��D�8�/�W���6��x��b��:��g�;X曒� (��+w�}���lu��+Pɢ���+��]��,�?{#�����Y�h�����շ�7N�m<�l�e�EȄL�yP�C8"��w A�@>�~�U!�Y��jEՂ�%��*��$7'�)��!�N��y?����(a��a�_<S�4A:�^\VT�D̘"�Ne�Eߕ2�]ϟ��({������A���*����K/�B�3��uYB�ҫ�i 5�TGA���6B�I0���_�N� v�kԑ�07��"�љ��\�87����lE���jVR�z� �z	��� }/p0�a�T�s�KU_�Ϳ��Q ?;�*�#����u��Ec,����Sf���GI��:��E p��!�3����W�R�?޽��[yqϩ_-,�{T���&��}]1����4I�l`J�үm��m��k�z�Â(��q�V�L�%��ݖ0[���q�h�Y�Yʧ��K�{s��=����L��+�' R^jvr�qy fC���o��\1|x�T"H޷��;T�_�B{� �����W�����^�(�`����!�`H;��Uf� &�r�<B�I� �*Ci�o6@��Ǽ�߳��5��n	�H5?'��o�������(:�0;�E�i����':�ߝjm�Z��Wh�
�����i`�q��y~�cc���~N�)\3`�����7/>��3�~�GY����wg��O�����\�J��*17zM�h����Dmꋻ������k�{h��׹�Jˑ��<���0��I���o��ص�ʗ/u�FBN;ÒÞ9����Կ>vv��U�q��T��e�����c��^p�"��u���	;~&��+�dP0�.�펴]�Xފ��ދ����u6�"��G�0�a5 ���36��[�k͆��-��W7RuH�^:K�hُhR1�!�g��`�{(<���Q���|f���� Ņ�!K`�w�٫.�H=j�|$ع�Kt	�F�������n�K�� ���d"R(��=I�;�zΙ����a�)�΃M�r�2J^7�J���,6��.Y�����)U�mHo�5�N� �,W�l�^��1�NG��������1qz��!	�&~���39�_Ȼf���!a�W���v��I޾0\�>.�P`?���'��Y�]��c<+����\9�u��C��j��c.k�4_�
\o��@�m�7�Lz�P�8*#/	�/J,��P�C���h
����7�TW�*�˦��wIi����wS`�_��� ��#D���NU��K�2ӊ2�鯚15��i���s���w�f��8� ��ƌ��]Y�ؖ����$yl47�R,��9�X�z��H;:&�4���˯��̾��?a(�����[���/��,�qzZ�O�Oz�N,'��O$X�G�w�,*B�`����SQ��΁C'8{�L��@	���K x0?�U�,�� P�w� �]����O���lG~�v�-�޷�|<�R�16/A��ع���D!A8�0�o/��JZ>#�0�emN�@v�g6{���c�QMc��$�7}(�1�P�ZUK=�����y+n}�'���*��5�pB�f|�5{���|�����;2t�嗸Q�c	bE����e�"$�]�?�w�>xk6e��ط�� ��X7k+��1����'������i6���E��m���π������������O}+���M�2[�ԦO�>ȟpq||zo@S�9�]7����קq>2�u) ���&摇�J�lֹ1Z�g��R
8#@a	Z���ѱ��W��2��<3Pz�`�DUC��`r�� \���A�I� ��&,�,=j��P���g�z�_��)��t��*����K�����O-x��Y*X
�-'9 !��O04fD�V%T��c׫&�A��]Y������Y:~���З�2v
f	kd���%��yt��������=;�V��Ja�	��Hӕ-��$�~,@z�%A���{��� �-d�AŎ�ӑ��J��6�m]s��;���uf͒��Hp?��6܀��y-P:�JG�g�3�}9k����[柮�x�-�0;,U�ъi%�ß�0Q����X�>�`跌%P�q��[|;T*���_�s� �t��A2&�0��c��o��|��b��g�L�u;��K�z9 Sh�ZK�)�	���J��%:6��[��*@���7�-�����S���׍<�n*��4�_����+΢<:�p���ә���ˌ� �=t�Z�^ih��:L���KW9d����S�Pm�����Ǔ�O���썙�4�����3�Tե�mb�s����ie���~]��G�Ɂ @�r���Vi��h�c��ܨ�f�"6{�*�6��OZ7�?w��̐-�!�yB,5�2*��p��Q��3��A0���XM��Q�^˒*jQ
1b�K� !� %�?h�3Y��}�<�41��­c�4����v������{�/#����B�'�Q�.��|�ؙ��jh�b�9�'s�/�L��.�6K�Ո{�̑ ����؛w(�Tf.�\�L�.,���V�
o�6�=Ss �����ˮtF�����p�bdZ��1kh�z8=>��W{��L=}*�uM�F'�p�@]����T�6��1�Lt�^�����<+�@�����#G �?ϐ�v�nR���>\7#��4�[���T'�Z�.�%ס1/	��Ƅq>PWw�U���[�ض5[ͳ��@��ޏ��s<�J���]���:0�\}����)�\��W��<pU����k.�^G+͢�p S4��D���a5�Hj$�� �T2͵d��9���=/9c	�b����y���i�J�w��v����x*�ģ�F@���X):vh�^�S�dBy��$6L+}�*��s!s����`��S��jBa�R���4&*V�&v��vS���%���4�}׶A��C��z����;D�<��x!��|�?�,��0�H��tK�X��H�5Z���q���T�o�ڿ5��-� P@� ~Hˈ�ⓕ�@� �5�m�4^<|SpF��qB&��
���ݩ�uLa��_F9o�XNwW��ϝ�F��T<�$��s.�����9Z���)Ks5�q�>5*�M�������]���k�y離�� �j�x|�@uǠ5�$rh�F=��4���T����4�ZA����-*'�ʓ(}Y���i�`�?DS���l�+ٙ��d��U,�(��H1a����a�4ʐ�U�ĥMg��qYK�����37o�6��}��ֿ{&M��O���[��Qo�W|MX����z���2��.��V�b��ݽ��b�S�,�=V55�CY�����D+�6/%��b�?��K�[��9|���%H�]�a�������kPc�Z���C������0#���5�f_�䜑l��8����q����ψiw �q��H��ga����IoU�8�p=�}�U�v�]87����]��:�y^VV��U����ۮ2�4ڤ+^Fa��� �
��Q/�$-h�#|�<�}������FV!�K�j<�;��
_Wn��v������(Ym�5f��(�v�9�����K�utЦI���ߪ7��%����?ai3�����G��Eg�2�r"���JF���)��,y��; xS�!_#f1�/�L�F(��*װ�ksAL^,0�՘Q�>a ��ˬ�+�M#���ߩ��\�H6E�1z- 4�E]��Ө8�吐�s0r�R�L@�< ����c?B	\v��gY�2sy�n����#��F���t?}�R$�tp�	�/V���$N?��C�v�EԇzZL/�aT�@؈',a��U�牕�v=�öv�/�g� r�f�J<x�&X���es3r�3��Y��;�����w{n�-6�e����XC5��P�����e�9��*�R?=�f���� �1��O��c?���B,M�N0��C�&���)��`W��,��w��E�N��ުJXUߣ\pYr�UGV1bg8-�SڽkE`$�AZ:[Qj�u���N9��Y�6?�L�'�'A��qSVB���K_�=ܰ��_�!V]'G3�1�H���I�+S:w�M6o��<�Dwr�*aY�X����s"�*Hmjp�WZ�\D����BoNHL'W���i�+�L�gN �����Ve�i�͘���픀�N���3b�D�-��-� �)��Q�3��^��s���Y�g�q*L��
L��M���t��nI���B٦�z]��z���ȩ�ҥl��+`�f�w�$��f�/q���ꂒ;C(������}�ѽ��*�1�cY�C���a���c��)�Ϳ��Pe�Ԑۚ}f\�`���р��0��1��V�X�L<�'��E�Ӫب.G�	Ҁ��A����$�0�k:gS�%�M�`\wQ�U&�h�e0F���nE�5�e�ܤv
��A��_~m��/S�Z
�U/��q��F�[:\�OD�����V������l�QO�5<��+���2�D�Q����խ�������EV^p_��V�g�c	R58�d��Ǽ�Y�=���[#$S�^���y�&�2���4ma	w����	DǠ{W��TI_	�z���n3�Z��}�d)��w�[������>����$���lW��9 �a$C��o|B樍h"�U�ҎJ2-�m����h�!Q��}q�1
Q��3M�=Xےk���|b�uO������ӑ�ظ�΅�6<������q|��gʹ��b7��w��ˌ��.��j�'t�}�����,'�+H�&DP�U�����N� ��>ϭJ�'pv��'�cFg����,~�)��u p��n&<nf��HA�'�:k�7��u<�_%�Gty7w�����0C���+{U����z��Km����K�if�^�>�����:��}�޴,ϊh�Dy	g�8W
��ʢ��S���o�Qy:���EQz{z��͖�N�M�\=~Ƙ�g��\�2�	u4������}��b���v��Ji���!K�]�\j˨P:��|H7�ĩ0R��x6���#s^�J��,J����u�,�D׍M�Qv��tb�s/�4��冋O23�b�������a�P�
��.��4Pw��6]��0�P���'����c���n0�P��4�/�9���U����"<��8����"X�z�6��$��i���4�Npe�	e�$����2���V�Q�RM�n����� t�O����'�!��C�m�/��=x
5��޼��h�}�3*�"xp�{����C�:0|��M!� M,��,��*���R����l�ݸ��ՠ�w��0��Uh
�.�,Y���L���UGR�h�W8���y%j��"���W-�2��QAFx��g��zA�dO�g����ɫY#����%�H,�8w��߱��,CW�����l;�מ��V�A����U[u�1���+#���� ���6�����!+�0�,�����Z�gr���P�du�
)��އZ\k*��鹤�׍
4.���z��=��Pe�&�؊�:K�}�[/�e�yo)@>UW+79ȁ�U�T����@�f�������y����t��;Ud�%�͞c����<�G��
��BK���H_w�k<�~�Y��]�v~��M�#I��W�#m5/���y�4�V���V(9�~�1��lP�$��6E��0��Ě�Qά�͆*=�OLUa�x�3��g���8V@��'�􎴩BX��w��Q5*N�?���=_�������lK�.~�R<�HN^�IM�����m��!�����N#�2cX����ðf�G"ոP���9iZR��n���j�V�w4��h
���U�ɀ �J^�!*a��c���Bb�+U������:�7��ʨ�:ͪ������bQ��^i�D�9�37lR�#�D��Y��xjY�>�&l�Ȁ6T�yq�l��l�~a��=���Y+]<�
���O��ʮ�7}���~���Ҟ�����o,�c�0�e5���R���\*��%��I��&�#?׈Dh���C���H�	p��<f��<��I���Fd�#Jt��*E��a��Ӆ�Zg��=�J��<��5�%G`B��|syx�?�޸W���	U�@����΋��ʜ��YHר�a�#�R�)?�܊[f��{��"�� <�����uv����p��h�s��=�d��:y
0���.�� ���:���k�9v�����'u��2o;�e}\�*���M�B�HlõUi��?��cp��M���aK�g!���0G�㝰�3�e�2]/�hM11�(��L��<K���[�Ո|��'�Z��x*a�*;�^�r�[�����^F<��� ct�5��pI�qS�!$�������8�4K(���R���f��6L�h ����������X<أ؁�u+�ɮ �L�=q��x�����٢C���tK��+�����V��fz�����(��#�q�F(�]�$���Eދ�Z?8ǝ��]� P�M�܈.�H��BNjT��XA�1�fJQ��^̻r�"���c�.������s�ٔ��f]U@��a�|:�!�Z�Iӫ�so�ղ��ג��oo �qIY��7
�*�%��L+P}0�j`�0�V�Z����<�W���@w�lpb�Ѱ���%I-��fCfD��j���}�����GK�v��J�5��Ϝ+'x��������v����q�?Ҋ׭M�P�f��l�D��md.��m�$����<�t�˘�Q����^^���dW���~%YjL$tR�]�ڂ<���kE^b�I,tk� �<�VC�+�Y�0���\6TЮ��,���o�fXأ+y���d8OQ���3���e�O�>�_�GP�v����(�}e���pkY�^?�61���x�N\JQP&0�;U����E�K�d�規 |)���e�vVI��hg�-��&DU�d�E$���0�A�i�b��+�v���L=��y�0�D���j�6�mF��͑�.�="I\��i���ǎ�1�����/.����=��A�$�?F��� �X~C�X ����+��)hz�����u�-����}��e�
ꇫJYB2��n�y���}�'��{�0�4ϱ��.��=���j�B���4mj3����ֆohj�P
�� 
� _� ��:��%.���r�H̱�
��\�\Y����}D9��Y�%'/1��9geF-�[�����Y�v~���$�+�/Ⱥ�8���4,f�sl����ϐ��k좃ww:G�A/��kȞ�P�mGt#Zu�Bҙ^[��y�jy������Y��Ώ�9k�׆�88���y�f.c�=Aۢg%z##��3Jj�(�w0p��5T��w�߃L}�F�X ��$�fҠB�g<��[��\
K#�-�J��׮	���6@���a� ��������М\rr�~�]K�қ�ދVR�4r6s��@_z`�p��`���C������W�mn��u��P���"�i�./��R ��	�	t������5�����f����H��Q�ԥ���E�;v;&]�rJ�Q�M�ž4�d�x��!}��(ED{�����h�4-�hc�Nʙs�Ϝ�X�K�g	ֺ�ĕ��1߉i"^O�n���{`lY�i<��Οo� �f͹���^�'6�4F����W���@��jR�p���<.�L��)���/'�;�U�]��Ȅ�1����xz�6#�F��Q\��w�̝cBN	il��<䆝|Τ�_�`t�¥�bK��n�ľ\hIP�V�$������A��F���U�ux��;��'U�@�b7`\n؋���;a͒���J2yH��/���Q
u����9��|��\����}�NN������%mr^��u�qx颰�9��\	u<(@�]*O<ã7,j�2҉;@G��aɛ����ʏ�C}f�H~���&����Cm�о^ͫ�4P8.����/����V�@|���Z	/V̻Z;IBfqw�wة�'�%�&���P�N$��a1r`��\�-�۞}Ⲃ�R��_Q�Ծ@��x�����Zd����O2t���rU",��lj+���9Б�;�TM�t�����rA>���c���:��.�����6ɵJ��r"�����l���'���3�^k�+h\�1�`TV&��,�Ju��?*�>
���~q���6iK	��}��|@�.k���7l��'�i�UXHM鱶�'�f*4��p���.L=w�n�����p�Y�o|�t�� �FP�"�	��E�n��I�|}]�!e��)C}�٪��U«bI����q�ʊ�t����_8`�q�9_q'm�Aa�6��Kw��q���R�T��5n�A�Ia^�rO�0��N������	v.�d�!< PP��0�}+��@�	���S�հ�A��q`D�\�F��k��'*���=>Qq�\6�>�����3���rdj�%�6�S���g����^G��K�f�������s/�8�2��̈�yŹ�K�H((�Xc��kz��z�6�f��Ϣ#�jZ��[�@н�>d��� &�Ds���qn��i��K#� KX�6,��Ȁ��7��D7�-����������I@��/N#X8ؗܒ�+������#%pp�8yY��]����S�]��� �����~T���,�2��s��0{��|����1��7��:�O����&�h��b�S�������p����f���D��h{T*Ϯ��B\��W�����#Ւ'�!��At�QdRK���`udfA�B|���g����nߥMxa��-I]uK��L��W�Ϲ�V����<&�@+mCO�#�/��K��[� �:a���:Cx!�ѫkZ����TVR	��Nݳ�z���1���<K����1'�=��6���=�$��ɨ��傓��V��
?��o�)���Pc���L@�[�r��>t�I#���P�<7�����BO�� M�$eo�2)qlZ�)|!�V�h�v��6]����磁#I�_��6�[��q�sAe�J'$�hU+
Ј���.���:��?bФ*�Oy��Ua��5+K�tyg*8���O>	y7L<�M9���L"�7������x��T��O=�biW���p8P��ގ�7�I?�|n���$�?i��>����8@*'�\�`��0d��F�[S�L�{�ΛƂx�&�e$��c�N�o~n^�S�[�&��#va�Y�Q�ƌ��{�P��	�Uq�~ơ�����[������s�VIo7��#��b�/���)آ`��>.������	��k���t�K��������@�ZI>�%�l~��"��8���BJ� ��Bieہx�l6CF�V���N�����{�Xͧ�V�mG�����M��#.T(��:��$�OEoM%(8������ͼ��IA�a����aQ�)1�U��T���z[�&t�z�:�${���^���G�	YV�R�CzN�F��70q:� �Z�
y��i�Υig�|M��FB��3:&ؑ��ߡ�P�ª������
r/0Y��c���ӎ���q*`���֎�Gf6U�y�5���G%��!�?�Ea͆�io����q�����v�S>�E����kTu|�B��"��	��J['�c��|��$l�a¥C� ��瞘K1�Jfw"r�
�]�t6�hC��'<`�qZ{,A/�)\� f��9v^X*q+2a�<_�F�΄e����?�U�P&I�gO������4;yJ����̰�8����l��1Ζ�]?����ٖ��;.����Y
X8�#���8E�"� q��N��ƎX�2��6.T�Ah���UlE���b�E�˥���z'��f^�3�|�H4��`r1�h�θ�c?��|�㢵�����:,�lYW�Α��,�U�ˈV�|�/,��yc1�ֽ^��|�C��h�́�\�;�y�qE����^�
^<�UԈ �ò�L���M8�t�f4ݽ�L���	��x��v��,vf�t��98�X����Ɇ�h��B�ӗ��0)�tK �����z�.��+nGt"EE�{� �,��Xi�Z�Qc�c.!m�Y��ϼ�t��Ys�>*V�k.f�ed[�37=����پ�J.��R�1��t�ݿ��_4)ֱڠ`���?�F��!��
��D�����x�6~�������|Eߠ�2�(kw�!G���oYխcO&2��*�w�p+�q���-T��ڎ�l���qO$��zY\�Xxi�)Y�y���ƍ�lS��o_`��3[��஢��a��J��/y�0r)]	��2W-̫��w4��BEIsC���j��龽�P�o�N.�IBc�k��;S���R��� z��9��e)��U�ʻQ�4A����I,I?]3�㨠�ئé�=�y�8�1�9����Mj!!r�EE���8݅�a
�w�4��M�_�{;h` WV�v"z���Y�RJ����Er�S��Q���$bh�2L�ދ�crq��U
K�A�q��o���E���ބ)��T0�]g��Aׄ��U�id����G�s�4���[/Q��Pa�eBao[�������~m�$엂)]��MJ�s�����ħo)���S�r-�j��fU?8H�!(�ם(@c軬'j�$�=���8֧�M�)ç�Ë@�i���^1~�]�𽰔l�r�6�+�JT�P���w��@A/F����ʓd�UOK�)��+���N��qW�>��I���W�wc�1��aF����ˇ�s[Д(s�}_޺xʈ��^>e}����u=���w���V�/���.K����A���<�x5
��p�� �����Z[ʤY3R:��Uq�꧄lX������(��xY�<(T,ѡ����BQRq���=t�K��%�uf�D��ɩ�xX�q�*�Ğ�Y�œ`��$o�^E,a;2O2E�{�R[d�8u�
E����P-< )$���8=�pk����2_��n�P�j��F_<ma�H=�$��z�k(��r��ѨǶ��Eu;����`PBaKR���yR�>�P�/)=��g�j�<��L"���&��%v�������!!ב���N5�w��Sj��4��݈�d���
ohS
.^����n���-�h���|�0��t�X��B�������g�);Ţ��Y6�ն�>`��[3�_�%wH�rS�����#_�u5�X��f�A�;��*�`�W�����&�6G������� �E�9��+`�x.9���$T�*�����9�4�Pf�6)�}k��xߖgS/q��.XN]��Gﮠ��������p��>�jı��2/r��*/,��O�F��;<�7v��ȟ�1>�ʁ�U[Xk���#�S]e��$T��wމ�h��
1�H�`	�b�J����4��`�\-��b|[ŏ��SZ�\DvSYu�.a��Q֒u�	g����9"A�v��~D��u�@���͂ŻG\�_1'�:�z�@���Ġ�.�Fp��rs�K
\5��,�f�J�\p�ʨ:�0"���庰����c��ƭ'a�{<�{}�(Y	���4c��
/Kb�fC�m�\�w�
�ղآJ;&�
]�!Mu �����[��((�9�	�OXG5��(i8i���ܕ�'}��;���4h���>4&RN��W��.� R��3�5��h���"���G�ea�f�N/.��>�(~N7I悱/
Py�M&�Ev&��=DR*}B��s��������˘4a�
����z����x����#����=�Ԧ�a#�L��.B��&Mp�IŹ��3�ì(��W��)�����\����~�I��j"���q&���#�V��?[9�'�xM�R�6+�ts�h�+��\������g�0 B�W�X�"@���������ʡ`�C[�׊Ց�z�<�v!`���P���Hw&Q\�(�[DI�+�Nf�Y�4P~��
2L�2�6Yߤ��=��� Q
�4�pz�'&;å�2o&+c��,�z*�7�1�5��}���`q�4@���굆�ih��4柙[|��!�<�!���Ѹz�8�5upA���BC�e38B��/Һ��A�ǉ�s�uf�""�Nm�J�B�� �u`�_�$� ��l�0�*��?���v�:��?=���a�f9���1��Ԭ�=
h�#�{����EJ�rj;?��`-�X�T��l��l`<`|� P�BZ�p����Bxf����D�[��@ya��h�"�W��6�?C�XǍ��4�l\kg*Co�����EL�j|8.;.B:���S���%O��%lA��/|�q��J��h��wZ������ �Q&�E���A�VTQ�+Y�]'q�a.)���`~+�Ad'��Z����Z���&v@�����(h|�&h3����e���,5ϖ�Bf�1���ɡXg�.M�2h�\#�����i\s�����m2x��3��,���L0��|E���o��;+np����!*�ų{%��$3��ol��0�@�gpZ���+��o�`Iz卸8�� a,x�vO&�е.�HLVs"�-�䘸!4�~�V����&�"<�1|Л�ڶP��{l�Ch����F�ood�ģ���pU@I9�D�ΐm�3р���39P�j���+�Q�q�!�Qg':a*��Px��l�Ac�X���.�gXi�`N�o�#�ZrC٨s5>g��2�
���{$��1�r�a��c"�ۿ��y����'�B��:$�����Q�87��%v����|�k��g^ J��>�`� J>�G���Y2��}	a��L�ξ�V�ɖqN=Ɓ�����
h������s��so���tC���xN��i�\�ָM��cz�$L���|� ��L�5�i�T�)#� 8�Y���xA����v�ϥ�$�������O�`�S�}�|=xA�r�5�鄉���#O,��n �.*H9�6�&�{6n��U�{$�>��K�4�O?0�/�ևM�w��s���7P��f[0�[Yՙ|��L
OS�g"�}�!Ć`mZ����V����(T��Bn�K��\�EN��d�?��0:ԑ�����R��/7��5ɘ�ֻGI6�|���8�Ĝ{|ׂu���H�x�9�zǍ��,�CG�^�F̎Ҙ>F1\`W�O�p�Xe��oY.`��(�d�w�����eXf��󉛇��tH�%He-;��ղ�tu':+H�� ��׽��~!�ؼJ����e�[RmyE*�YW���?~�=&,ⱖ��y_���ޮj��b�X��J�ֳ�叭"����gf��d��vÚ�sa�x�d�U.�$U�u||�{�i�Rǖ���������И�g�2.���߾:�4*�4�
|
��C���=2{z��
ݤ�.����dv�UXK�9�� \�3y�CP��I�jb����G�CU��Ys�Q���	cV��JY�6�����WY���C۾D���k�}�o5��[�s��g�g[όZߜ\�h�x��z���(�~��h�����=�ƃK����73�7����L�T�3��Ǉ(��yem@�_]��bX�j��n a5Yϸ:����V��p_�
qi8��@1�\�U�Xz���tf���tZ�B����{�l&�`@�`��b����nuߍxFϺ-<�����h�<�A.���J����7}i�a�N̓�q�Z)��n2�c��l���>�1w�h��jm�ɟg��x֨
�.�WFǙS�0\��T0#���W�3ޓ��,�C��Kh��CUC@+-�և ���\���ߑ}���שñf�?�^�Ȍ{l�p���-���}��M����%ؑ���R�n+��>tEۀ�6\�����^l�al�F7ˆۊ�w��������tr�Hu��v�/˯Г�2(׳�F�{�_Q�uGt����y��8)�)b�F-���iץ�^�O�S\��du���J�zrW�
	h�}k�0N�.m�9�Dl�gG(Qz���F��A�N5gP��^��*��t�G��2�v��Q��3H��@#�H���&j��Ί~��p���y�30�a��~<���K�j�VԿ�~���[�������D6�4�C�+��Jnp�����j�X�s���V�,R��]�I�V���?���AL/U(wZ�cX�B'�4N;>4V}�?9ы�6���mR��Z�|�Q�L�������.tc�kthu��*5��mr�sڶ��(AM�o�qo����O��"�rܘL}�]W�AЦ�q�	��25���
�\ b��X5m��I-��DI���� ;�(Ry�����RvC��`�zA.����\0>ѣX �Pl�\.��atr��%^������cj�Sq�7O�	_�D^������t������G�E�KX%&�Eyw��s���|�IB�5�7_�t<��Y��Œl tF����&S��2���W_2ꯏ,�ETȐ����d�
j
���k��Ȓ�a"��L]�+Z���2���" �щ�i������D=��^n��]]XD�����-���f��{� (ҥ[i�N��?$�n�e��U�]�L8����Rnmw��G��ie�y����G�nW'��!<b��9�^��Z.#�o'�*}#���Pm']���/IM,���#�"���E���Y�����4�>�dم�NO���<�4�#|�~���3|��^��H`CV�Æ@%����/"��0��T�ʡ�V�%�8b�H���������������a4��ex�z;�b�^au@z��&�@����"5�vP"��*��[���p��K��z"�-�LY�|��s��1ow9f��f��ay��3!��W���b����>is��m|K<?��5=n$� Q��&cp�^���ad3��C�g��<bo��76�N�.�F�)��2�T"κ�9�t�+v��"�֘3o�H��z@���*w[ؓ�l�QTk�,��;��7xFv��Nm���Y��ԜM�k#�M���c�ON6ZQ�@����;�2>���i��R��eԎ��x�*��Nؽ�y��jE����FO��o�;-���J�.vآD'q0�ł?���_Ģ�iQ�[g"fd[���d�zVn����D�|f�@�nm��|7�btv��Q����,d���?��$����'Y��c����@����	�7�Q�*@.�W&��%��_x���/�^V �J��9�y_ٵ�����vk�
����}�Yz\0�}�[gZ�<�p28ԏ��5	8��9��DU1����Ȟ�X��#F��3������O�������Y�
�d,��t�O	��I芆Bt�vj(L�N5�-zb�R6�邿�Pa\_8,}Q�P���9͵HP{�i'
�m6�3�yEU!|� �
�*���l�M��7�[WƑ1X����P�����Ì��0i����j�MD����8jzv:槶}�<�c��"i��
�_��6�Nv�f�̯Η0>E]4AQA��N�#`(�m��TP���5��88�vUQV��s�2�,z_�Ɓ�����F�u#L�z���}yB40���ĦN[倔D�ٞp��Se4��4�g}F�Y�Q�
�<W��$�pIaY,D"]a�,(�~��U���=fP	p���W+J�ʇ0�C�_/5G��V�. ������fhG���^���i�����z:�]��`C�����?G�m���ד��{1���ݼ;������~�%��j�Y�2H��  e���h=WQ����ܰF�{��3��s�P�j��LwD-���ml
{����F�P!1+�R7z`���e��3�Ӕ�'˯�xZ]LO}���{�b�.�͝�w�Q�������B��U��w4B�����%�vh��i1�Qj����dS�����b� �[�~��e�k��TjHu��Qy
��s�w���K�Wٜtt���K����#�x���E�k��}v�h�i�-%�kd����1�[H��0� �z�c7,EA[��e�7�����HYf�%���('h2�����@#2�Y�<�KP`4����"2�8�X�������ƫǁ���L�2�X�cL�=ݸ��;<N��ɄS2���K�NAME��J=a/��H��	��]�����\\k�`A�ӵ>���te���.V����J8p��l�^^�j7��j���#�l>$ �H-3�=�������Y�6A��o�Û.iģ��OG����d`��4��w�D����a�t>���NC,���Վ���\���`�.��X����Tc�
m�v��,_�(����r�ɽ��5��w��biQ�O~� f�C(=�Da�/�N���Ɉ�䅼ЈeԁF�Ўs�aj�py��O�w����&�ƚ����� E^��ƃ�h,�����Q,SFkS�Ե ���5}-gHP�[τ;C�ZA��8�xe�4{���_a_�RC����r���1h��?E"X�.�(?7�7gP��{��93%+/��FZqL.�@>�ά�C�ձ��SXuuf���w��/�LE:���m~��g�����{�g�}Oe��7ڇ����`Hp�(�^<paܣ${e�q�t��Ku�`Մ�����G/n9���n�+��m�Tq���	�y� =���>���(W���w5а폁Ϩ oI�d�A(�i�,+Z�l�:&���h�N/֏�{��"�,���E��dxzr��+2��;W�ڪ�����݋)��wc\�*�*����el7q��)�<�g�3l��\@���`���Χ����Lp�"(ԍ���<�?������ɉ����Z� �No��_�Ɏ�2\7��9�A���r���Ñ�MGϛ���������/�����	h��~Fo�eS�jѠ�i+���&XFv`�̙��uO��N�k�L��<`��Nqs����x���AẌ���9օJTI<-ї���>'Q!"�J�>�)�zd0���\���?�I�s���vޅzv%��7a�8~D>Е3o�q��8�u<�e_;<�5�{p���GoI$W��
��M��۠Ա�#"s���N?Zg^��{�0�o�c��E��d�7����o�99P���R�p�>C8��yiV�b䋖��Re�sf&�.F�ԿB��W�d�k������9�U޿3���Y�\(���;�S�������*00$�l�A^_�pď�oYq,���9̣�}>
k]j���	YPbK�"�n�}{�Z��[�,N��~�>����KxU��1F���튪`�ܞ��x呴�9*a:���)���:e5��<[���u����|��u"!W��zi�:RX���pP��")����pσ�	 ��sG�9��:�9JX}��C��\#�E�F����8F>�7�*�����S���P7"�i��g�.�/��a�2�,pC=��c(������s�g�&��݌��+J�{Mpo\�V��9SlJTJ��֙�6�f�b��k��q>4R?5�?�"�ӹ�@�7B�@�&�$	�u����U0O.EP%�_Z	��7 �&�ԵX����/@O('�L eY�	7"_:R��/�nI-�딐R{iM4��|0�z�3�������b{R�_���dz���l��/<���Z��N��	�(n��T4{��~>�}�d����gűi��9ͯ����U�$���W�/ӟ�b�'noZ���)���T�����Ub�i"fև7�����y{�B�@`OΖ�~a-��D7j��a����%�lڡ�6�Z�*.}1�|Gs���l`�Q��jЏ�0�Gz����ܔ ��TU��w��D�}7k�s�o�������ơ�ɑ�Ҋ!�h�Ǩ����T>���e��x�Ƙk��6#_�?GwKP�Ɨx�S���U8�d��K�MT3�l��x
�vڔC_�����r4������� �Я��4�ͪrs��^у�WI�E-�إ+[����Å3�_LI����'Ͳ���<,8��f���|Ļ�JA����y��r"�2�d����ر��u�Q[�:1N<�,���Ҫc$%�A0ë����\�~��S��H"������������_����3�f*>}�BX�g*�n�!z���?�����΁�
x1n*�e��c��%֊r� :nR"	�l
�tӲ�}��@�X\j���4G��Y�̜��0�7��ן�8�^�_M����}g=~���fe/ǧ�o�%o�'�Br���S���A���@�Ț��N(��b�X�}�3��xc#.aL�z{��I0�v��PxȯQA�rwH�P2���?��B�lQ42؆'�:�.��A��5�Xm������J��6/D�תƽ8��5	(WLyj�m��m/m?&��4��^�o��X �܂�̌��ݢ�>p��mk)l#M�K� �Np�f�?p��^,��.x�SX�A�������$��վ#%��>�N��0�,��ˢ��7�I4��b�$s!���g�[����+��3~So����e�P�ƒ�R�	8����Q����퇅�PTT\��jFN���t��3��rF�]f�X�v������Fq�}����CdE��}�HC]6�'a��5T_3�5h��S���տ�@L�-w����|AxaE�7C���=(	��X2��վ���������\u�,"[�-��ύ!�b�������Zu��XA������ܽӏ��4T�����c��3�|��zhmn�)�&W
Ư�O���ng�V)3�+�IX����B)~Th�Q:*O��W�z����H&5�L�`�6;yz�g�5�+m���7���Eސ�>5cxn/�}7Դ�잲/����\NJ�a�WP{=\g�gi�w�`e`n�h��^��`[�\..P:T�% ���*�37�b8��N�\ss/��`Fd#�1Pn�m���C���ǟ�[:�D��j�ͼ��Qb>K;��K#E�޿��j����<
L}��=Hfj�3�8"�R��:)϶(B"���d���%���[eB����H������+>��b�,]���1^��㴿��5��`���]�(�'ch�cm`���-�|4~9CY��<���o�b�^�u�ז�t�pp��ȭUΥ�f�ݩp��}C(�,���N�V+�����<�s�/��!��8�H���~k���$:7�6�Ȍ�Ȣ ��!�%�yR�yy�ޅiҜ�����z���*�	���.��@��#cX�� ��ｃ����A=<)�!�-^���aQ2;��"ϟ��@I`�)�a�>ܷ��o�a�`��U�w���F!-?�UP�)�q�|W��śV�q) �"a��֋�=�2�y9�Yb�Bσ
�0ct�Tq�ݯ@���T3���Le�5�=��s �e�������fo�r�%�n�UX1�t>����Iu$ �Z�!D�Ǣu�>��H�G�Ut�_�o!$*9���ܴJ�ֿ.�)��؊Q���t�S�G=��@��:���dǓ^2�gr�F�4�Q�?��b�h柨@��K���sW��]?��D��Z����As�������7�Ŵ��$�I�T��y�>M�"�z�5"�X��]W�7��؝�w�[�P�3�`Z�6��QV+p�5�|���uJt��I,���|f^�8��+����O �u�c݊'�� ���8j`yU��l�[#�c��"�,�]���?l�mv'��P�Ǘa�����1H�SC#� ]�'�h�/'Ҝ�������B|��$�����0ya�h�v���Q_5����"ү7:3�s��e盡F��23���[e�&#j�*��;t��&��AR��ě�Y�>j:~%[��GK��d� e��_�?5��rJ��P�FEa�����៧�Qj��rp��{�xu,��!����W�`ͮvs��hJ�#�j��u:$\���6�ֆ��UƏ���t䲍�5E������Y�c�d)Ė3nKi`ђ��C�����+�hͧN�����H��_:��Rݍ��f�8q/����� a	зl�p�Ͻ���e�gXp�.��?W�1+|)ϊTk��:6C��
%-*�Ceb:��~����w��K�Ҳ� ���qI1d��Of\�F�������<Aް��N��Y�=ńFt��	�U�{�ʜ�7�Ƭ�R8��{ԥ�����F�6�����B\���蕳���K(�$��k�r��"E�f�G��\ ^���];�Jz�Hatg�ѯ2Y4��� A��o�{� ��C�W��y�~Q�sb�L��Q�1�1G[�$�p͐�	�����s� KV~OIi�zT��˧�$�n��\�V����E��"��a�#����C���z}-���5%)�)RD��n�Gd\�R%���i|flzߣ�F7�G���ߪl��N
�DŐB{�[��Ü�+W��@=���-�<���S��<��Q��S�[��$j�h���,!*��1��``�i����r����;]<hǅ�I�d�"3\�MS���2?�,��g��h���ȔC�ȶ"�b���.F�g�<��r�r&�p�{0��x����/�>�K�6�1��Y�í�*xy�����'�M�����~v�s���ٮy��l��� $�����1t�Ai� �1q�r�Qm��*�Z�C�D��2z�|���?~I���y�~���N2ѐwd-
t�E!l�:�J8�i?u���\��G|� p/lb=�6�ŷ��|t�4�h�N m�`gw��y�.>m�/_��D��H*'�����V���g�l~\8C�p�2t�g.���3�U�M']TM:�����L�l�Nh�!��~�;�Z���D�£қ�sz$,|e�ᬫn^1�,�b)� �ZM�;�Ř�����Ag��ǋ���C��g�l<+�eF�(�"y�V<�����)���5�J�0�
%��/Nt�F�����a]�U61؈��~�������ì9$��tжw�\y�4������[%f�ooT�S�u�+�GOF3M)��yL3�r"B���̛9��d3�D��3.4:Hq��/���>E<V7V��a�i���'m^�������V>�S� b?�|���#Y��^!.9�s�ؘ��#��b�)�I�`$�5�Gt�Ӆw1�s�u��\�w�̽�U���8���͡��z
Th���P�j�r�*�φ��zYQ����g��Kt�Ǒ�؞Z[�k[5��d��跢����rJ�ņ�Pϸ|��i��-��e�z-=� ��b]�D_�Y]+M�<��P9&���*��.|�"�M=��U43�72iON�ZA-���r���h<٭1��6˫���!"6�A��<yܲx��&�m�V�}�^�5���z}��
Z�+d�o�#���֮�1hS����g=?qf�O󸟍�Z��w]v~�y���H��l{-	e���0�C��p�_�uą��Tz��U��s�P�`񵓵m�ֳ�>�KA6��Hi�Ӓ,�
(�.N���q�(ǡ�T��y���4�9�guPŝ�
9�}�w��ᮬ�YjF��A[��m
Jw6*�G�P3rsr����\:�'��cW3Ǜkq�iB�4��͍��W}20��g���o��JnSR�sռ�%~�MV>U�q�\8��	�QX�����f����gq�#�f+�Z?����y+�f4dA�I����XuRq,'�AјP}��Sa$}� C�|��w�^��� �z�����P�
�j���8�Z	�Z�K����2���|����:�I�#1�ևm����z��|����o���7���h��c��#1��9 �����zV�Ҭ��!�����0����pX��Bk�N���-�� P�V��\ղ8۰جu��h�n��ĳ�a���B�w��nD3W�_�T�*��<�Eq6��{Ą�@�v.Eg~��T�м��VwV.Os�P��Fl�lcj����1
���o-T6q�g���5M�$x����A�ڙ�� ��7���k�BDi6	�l��?j��R��e�Pa%)�\���8��;bw��� )p�Bw��X�+zP�����ý���[��n�Z��;L8��
����pzƫ�@��O�ڬf�R��u�T�Z��f�F�I���vr���Fۃ>�#��ޔ��d��W]o�� `6t-���"N�|ϕ��Km��b@�yL�l���/��*�`��Z"&�Pфh�W�-\��_�7X�E�j����n����8���b�,?lgJ�GEB�Ь����V��:�)����C/�+���w<e�]����M ��lHD�$��S�	�%�*2꟧Q�Β&��*D��˂c��	��_�����?��+Bs��I���H`s{�n�R�gA�t�$�e��ύN�ô繶C)�#O���y�Л��	2.lٍ}jOu�J����9E]]ņ�~���Md(d^w��'deg^���b�''���_~i���J *��^oM���U�0��\1b�m���5���%��E�6�(s�Oϑ,M��dz�r�"�Vgo���f�
FF�X����"z����*�I�}����Óg���s��܅I�W���AB�;����[���!�^�9G��k�ƾ=�L�=�ǥ��h3M�
)<8���t�r��>(��U�uK��j��ս�����l���Z���K�wˍ1�ÄG�D�(���,�����B�Sm&�n��+��<7+�8�� ��b�ӳ�7k9��7����v|�7N!Gist�YтV̼N+��I�,E���ʘY�}&��o���D�5Dc��?>W�㷔�F{1��?6.��j�?h-����u6{��ڧ�0�v:ςţ@ǟ���b�4X�8������]��Q���H(�|��Ǝ0�Wg�w4�tD��A����M���+��U�kp�I�����N��a���N�^0Of�6Z-I���^, �U�1��D��k�v)<�D�"��������ח�2�2��T$��m�x� �����l�H4���>W�&��%K9��R2�Y)���HZ
�
m��?�?Vx�u���`�*D������s�����A�`�'t��{�Џ�P���뱜�(�R��+�ߵ�.Q�����al�d�i�G�<s�"<��}�?&�D��-����
2�r�,or�X�ŝ���W���̙��Wޥ[ZSao�Lt�4�4�7���w��`�GyW@��]w��xn�P�=߀��qw���Hj��9�=��OO�ˮ�Q|n���@�(t�#�P��� B�c�o��FQ�
ds�hU��S��5L��:�g�m�!P �?������pogC��ĝU�@�.။���t���+~�D���,Ӳ��A�J ,�f�d�]��	hK��9Z�� ���KN0+G��i�,�bL����Z���62�;�� �ݝ�<K,i��dQn�v{7���g�ȃ�&��n"�~�0@�TK�4KJr�� ʆݼę���ڂ�G�q�ct�����`%�w ��]��i�{�t���b�_F���wI��|Ĵ�F�L�:uAS5�C	�g� �7��Z&�#2e��1eA���z��V��\����E�J4��3W2l�E�`�:װ��N�S�^?o��icj4oG�SEVTF�3I�i7g�٧s� Ӭ�2/qE�s@�PR���l�N��Axn(���֍��I�K�h2���h$����s�1��߄.�3��e�L4��P����`E:����j���[�ݻ�A�s�ZN����Ie��n�y]j�D��Q���j�����䢒j�i�u�������U�TZSj�l�a�KI�����F�st)���K0v
�\'�w#������?�D1`{*�\ו[�6�sg�DX�}�@k��P��x^)��*��t��#�J�/��6P;`maŧ:@l�V� `�3�}�Wu2�xf�t�
����id����V�,� ���C�(����h�RoP��Fs�z�h`z=��%�$c��{�@�BG@� }���	8[���UCU��l�*��(���~N��Pր�/� tSr��.�G�]ҁh�
��r�Au������s�A6IPrO��7�5#�o 3��]uB�M�K�40���0��c��n^:��G$��X�j�sN�Z��ZF�Ӯǁq����n>����Ja+�Ry-������ŎǢ��O��v2�E�A����F�M���o=�Z?�8A�Z�-x�Z@u��z�ϙ2�uD���|4k*
{L�R&�n�G._6 C���i_�˿k&�e�~��"�>g���n[�L�{�&:|���r��j�{�@
�e�3�U������Y�~G����P��TB����B��s�H��m�=�Bz�2nP:8TeBݞ�|.��5%I$�td��6JN�=�Ɋe?7�o�����ᡩJۛK<ՋZ�c����:]�e��h�$Э��*xM��Կ��f�ˏ���̘ ^Xx�LG|*.W~���}����[�)}1ۡ��wa��S��	���6��l yn�6���G靵��b�$M=W��}'H>�ZY�
hO���j"l\ض�ǹJ��u��j�SpMiD��7�r�� v�8�v;jV��+ϳb7��4N�}����i�x)㘑K���z3`R�S��&��F�b�P�J_fN�^\�?�ܺ7lN�%�P�1\A?c��1�Fy]V�����oS^V��"ƴ,q��D��@� ��Fʲ����l��s"{%7pR|��_P��;T�c���'r��>&�4-ÁH�НݪO羢�{���xb����)���z*N
�U�z������@�oI�����`Y��5?TQr{h����Gz� ��U�5XH-]g�}�9�]R��K��~M,��^"Vפ9+זqD63���r���ט�󭸱���ؽ��m֐�����w7�vi�M�^��[w(G�.t�.�@�b��Y�e�>���P��&��l�������#'�}#^��1k� ˞o�I���,�i ʷ���:��ۓt����=BS˓�̽U��#,~�ܖ)�M���Ѳ��`�b�N����!t���A��A �!�I� 5���ʺ�\�?�;�7��1N�H�?IҞ@��ש��������Y�.��V�~�j�!	[$��v��2�Vv*2aHz-l'9�/�I�&�Ԉ� &h*a�G��@H��t�j��y`U�}0��'%���I�1Tvg�]d5���������K�L;�r�
8Yt}l�L�v��}�|Ex�����Ӌ�E1�ǾO8��w�T��8��]�q��m�j��~���}M�=�֖W�6+�%�P�{6��"3�D1��M �f�Y�����:�����L�����}
x��V�K�
c7���FI���V�w��ԑF�V=&YH7l����!(�P���$�TM����u����Q�_ͪ����vd����c�����j�����r��C������z�� "�ߒz��� ��;�K0=��<�
TQV̷b�I��n����4�o��Ђ���1��;>KKQf^@5uH�q��yuy*}C����C�ao�Ϛ>���(y�W���<1��&���K���e�.%�F�B�.}=��X���T-H3�!ͯs��WQ੤GM�k��L��>��m�_o���-��|_��+���MJZwO��U[0��k�B\�5�.���[�|���J�-���u�=��ۯx�P1�䜔)�n�j��~���&y��_)DowjJ	r�ct��`h|������1i�}�������toT�#)���(|,�M�W����%%�~%�]C(s��wBG��_F��]R"b�/�D�B;&3>���f�����NyX��9f���ư�Y�-�ĵ~]$�C��6k���1���%/�T�	���
�4g2���y�	0�3�m�;�v�t��Q�LX�rXQ��hr�ml����s� �`<������D@K����7�{ho��c���*��������ʿ	I��\�2׹�����J�8i�rh�V2��~���	��uᅈ/��qw$�}�
j׻��1�/F��0=���$�K���s3�`.�*X֟�M����A5���璝=e�����.�j�U�a���a$�z�c�IKͲ�?�KV��������B�~P���)f�z(t{���r��	��i[�ыx�>
���a�����?��pk�Kk¹���^���8���%�ʫz�[ɕ�C�e3�b�G@K��d���k~ES��J-l������!S��w`*1h���Ӥ�ŀx��q�w0��,W��0F��M|n\[,����Ԥy�QN8���R9������U��3"�6�j����y��Z@2A�ո�]U�$"ч�$}� P �
͠ ��&��`(̡��Er��7�%!��t��Ua6�K�&��<f�	"T��@]��R=V�+�|�;�g� �3{���7� Q.�W�Xȅ��I ����$S[�QA��m��{�6+�dD%�p�� ��O��+�\�M�e��U@���?U:ur��p��1���!a���32������*_q�
14���4�?/ż�@S��p,8��ϐ�-`ь{ciH��)�=�A�)����v�ʱ�õ߉��� &ؽWhF�W��DQ�������@g�:� u,��G���ˌ�5�\�&�Xu��|�������=n�OP�^����%+��STU�U{��L�#����w�_yh��9�s����~���PE�G��3v�-���B]-_5�ϒ�mQQtY�0�>���s�u@iZ&�/Ŋ!�f^z1��26�6N�=EƂPh�+���������'cF3�m�
�M�~t��4�.����R`q�Vz��bϧ�xԹ��&�'�bz�Zf�W��	���qϴ��� Q��r3�.�ёx<��b'_��a���L:oY���
���E
��W�����t$5�f-�5;�2�H��
�f��ZH<)is.�㕵%xJ*�ު�y�hՒ��-�f a���J����A׻�7#��}\?�B���"Uk2'���B��3�2��	e��T/M������![�٭��![����q��A��n�cI��u_���q�N���l3k����� �[��k��{�\���MIw�q�.����E�E��*BG���7�h]`C+��>���I��

� �Nxo� ��o��1k�b3T���Ֆ}�����O3q�Z��-،��b,�2$3��Q��8�b���,-�{ͅl�Й�{���I��X�Y����r�>6��Boǡߨ�8
 ë?2�:_�q��ݕ8�c�H��^�Ը�Xi/eJsU�8����ζ��e��y`��,���x�-I���<�r�b�0$��0�0���M�3��O�{�^���i�m��W����޳���C�،زVo?~\Y�4D�w�ؠ#��چ6�����~G4��ѯR� 7xB���Κ�<�(��՛�Q�����{(ȹ6��7���+���Y�HɅb%����5���s��Ֆ��忀n�n�W�M���]*�Y��i��(�|����������p���^����UC3娓C(���Av��]J�c�/��b�o�F���U �D��5l��;Z��Iw�>��1"Ġ<�p���|&i���Y�Q,d�$x��e�!� �ö"���*j̶�N�_Ĺ�0�_zD�]�����圊$0�rZ����l9���~�Kbs�+Ym����{5+�lcj�y�WF"�O�o@���_FO8D��x��⁆L� �ub8fHF��+����8�d�T�V~�v��;�����s��w��}��>��'�9���)!�!d�v�U#�/W�Kw���7�ּ!## ��UƏ�lɷ
$��W�k�:p�Y�u��f#�W\ؙ�8Z.��N,�5�_`4��?%C'-���5�����a<�{S��f�&F�)�j�V��ڌ&������{�2RY��	�f�Tc�Y�c1v�q��p�Gp�O��|��;���Lh���Y��"�?*�A�ԭ�liYHV�P�׉r�_v�{e����'��A�=�:;h��F'~��b�v�Zgۺ���|ާ�՛}��KE�)�=V��^0� a��r�da� ��\]��� ��Ukݭ�t�B��)�Ni��v�j�U3����(�@"$��y7&&�]c�n��ȶ�y��U�c��LK0f�ac7q�p%�c�dS5�}XO�[������dy��A?�F�ҿEA��'�hx�[����v`e4�r����v��3V��9�}`���I�en�8�^�}����)l!˻��Ϲ�.v�ݹ�|4`�mN$z�آw�~��B�q6lo[,����!�gZ�/����p}v E(�Q��I�9���֗��U��U�����	i:\��?~����C�^%�4�ex�*9�:(I��g4"�����Cy�^��@�ie�b���dO�\�$�a��	e�B�����c$�	�l6�8��\�W�$ 
؛/���4ж�r� '_wL�:|M���Fr�R=�#�d����5x�5�[E��\��8ͦ&�(ck؃�W\�ұ*�|o�7��Z&6$tx��'JY�\��>}�Ih�gTP��F���k��o"������i2E�y0#�&4��/�$���צ�㍪u�������qQ׋T��8�sU����@9�47^��4+$��dw���^�1]���)t�f&Z:Ɔ�e��b�S~V�g�����pHi�cPn� l�ڃɩ��,����o4�=���Hp����ʐՃ����#�ƶ} ���^��T�h��\��Tl�>sN<�]��߽d|�Ħ�=�����Ζ�H�����=��$E���R�D&&
f�����f���q?���'!�0<� �E�q�����>Ǣ��5����YQzuW��|��(�����@v7�.�a���ȋ<����/�q�7��q�6�J�:>�Dw�o�j�˶.��h�
\�}���l\Qt4+�ן�����닉�hˁB��"�5}N�^�Љ.�ca�/�by`�@���h��ݚ8uPo@�Ȑ3�̇7�P�mɶ��_#Z�@E�Nw����
ܮ��+U׊��]�3E�9�Ҍ�S�^7�`)����.��yyyT�$D��n�Fj�a�����.��cuɇě�����,�t;7�!Aŷ6�6�Ɩ�Zw�ۀ"����P!tʳp�ט�v�Rj����h�I$[�^D�]�3�)�Kjc�'���5RBd��"G�5���w�I;~DS���υ��=�BvSyj��$C��dؒ�X�wy����s)��E7�����xQg@��xO�-�H��5�L��gɿ���}�]�
#IE�s)m��GP�����p�N+�5��#�baK��0� ��qBpc�����K����u�؋�ȕFV*�-M�T�a�������T>`�1�J����� }�����1�2�5��ѷ�n$0��N����-�&��.��lZp�荾x������Ϳڪ�i"* ��2�6�
�gqJ��D�Ɉ�.���A;t�`�a��ԯc[���ٛ~�:[1�3��V�H���+)���!���5����������HP:F�%^7��m�t�+b޼$�:qcSBı�?K�v"*iU��N��#t}�d��t"yӮ��/!� *�`+�?ME A�WK��$��!G{]2��.��=XrkY���6��ڼ߾��ljo�(�&a&|�*
mT�L�9ul����sgP6�6W���&%�oB.ҌXd G^��q!���FƂ �� K��fo���+���K*]��p�&0��R�T�`��~��� V�
2�e
2�fR~�|7m� �4�͊�<��\Ŀ��^#�ξ˫�UTP����m���oB70@d�V!N�jsC�*�����bSS��U�"�7BRv?��i���c�b׵��K;�
l�3A,�K�nK)ꡝ&�rb�_bh��ʝ@w�\�b�;����Ģe)�y\���1035ȩR����b-�o_�`���HV1O�1���x)J�M�����8a����Iz&)r�lݢN��G��k�/^��"��㕟r��Ȋ�bűZ��<��`{连t���Jݵ�EM��
K +�2��c߈�X�b)��E�6�g��aU��3�e�D�0�[�ߘ��ax��˰�,��>�D~�x�{06i���l+�>�d�t���#��|��W'�.N��C	�i��oB�Z�/� z���!?i?qH���LN�έ>�|D��(q�u%fdrw\�OsH*�r�5]hYf%��cl�1�8�������.������Z����`�=�u�GԀ|�a	Q1�M��B���~J��m XO��ˁ����l����n̓ �;w�ҽu�/	JQR*K��D��sy
���]s��^ܳv�1��������uȅb��>l��
��3�W�Q|�~Yy7��4_�F�c�X+�Qgʦx�u|]p�F2A���;��}g�[��[ȅ�&<G��-=��� O*��^�176�+o����I��A�+�r��/�4�s�kW�=��U �������7�o���*��Ɣs�
�;�g&<��C��g\���w��R�<�H�~`%8��
��3��s���	flW��!D���6da�#��!W��{�<.^m�Pv����ΑTEr������}�B�I�^�41�|jdeZB��=Ю��$���)���𗰔ǅ����It�*��{8��m�IE��imt��X��~�+�.Fq��!}D�<s��,y��/f������+��3����;�\���UN�В�z2�l�����"�`D�ډ'�J$?�L(M��B)���k,���QA.�H���Tk�	ߎ,w)j|�Cw�y��$����>.$��{%����$:��{-���H���`��L�+�1��t#:B� 
'��ti�G>��F�q��)e }f���`�_�HD�؛+�݉Zô�cڳ�՗��Wa�����|�c^O���>��$�@��a�pwQ'���7����h�T�M�9�b~:�5�edQ��SօFQ.(��
&V�U;j�&��y<�o#,E�<M����[{̳u�!�P�y �
��q�̀ %Oj5��/����Ee�	��j��[�%���L�[ħ[�!ދ�gyq9����jyAW/y��D����t8���\>$���o��y���t����	%�T��n`�:�Sx��@�����8�x1"c�*�:��F:|ե�F_�*�mQ����aA��U���i:~[(�2_(
-�����d�����X�����(�ik%I���[lٺl��ٿ�s�U��ڥ��N���m�mH�i�G�,o���e&����,-��'ǩ�� ���K6'�^���1��Z)<)�y��I0��zHJ��P�x�er�u`�����pz/����B��~?	�tW���iPx�Gne#8�I"��>�c=V�T��|C�e� z�J�=@
ԙl<��-�s/%N�x}���.���������tTZp�ӫ���x�-��5#����ы��^��83���#��/�V&굊_��	\�3�iX�xdg4E��78T[�6�(1�x]�~�ZBO+}�3k��X�G�(�������O�(׆�]��'6!Z����fg�����
������xz�N�qNa��W����*q�]��xB�����Q�R����pM<f(Ѭ�3�%�}bO}w�9OYP��g?��l� `m�U ��@��æ�������Dp���Ƞ6W~V������  j�6I����}X�o��4��N�tv��
D�4� ���Q�hw�Y1�si2e~���! 8�Al�����c0me��\5{���1��%���zLR�� �k08�=]u��zWuLlה� ڄP�Q��k/Ď��i�⚞n��l~y#lܠ���n�G����Z�6*� �Z��ks+Zm�" �����	�J�-�iϊ
�/hC�}�"w��}��f��gܹ=ӕ��:�?�:�$<�|R��1GAʕ�{�7�.ڈKm�f�Z[�I���<��`�m#4=����P��vmweէ2$bpU$t��s�J?���Gd}�x�jJ86D�m��i�F<C��cV�~����Em��*�o��/=�V]��̚s�C��3����մ	6̔����,�,�L�0o�+h��~"�U@@5l��W_i,�>�841=�(��cDm�HR���L��_l?�*\ܳ[�K��WQ�l=�Z:ï}<�1��)��=��5�j�����LJ�טn�0� �1������K�wL�;�pH����-$��)+�Ӎ\�����\�X����+F\��&%�ek*v+��2��s`�a�p���w�+93N�S����@ %�M���#�A��e4i����D%�4�c��O�W���d���oY}�QB�?��$�ָ�ŮzN���)P)��o��@kyu&e~}1�oYlq��P���,���x�n�acӞy_V2Bb��������&������>3Ra�YT����.�d0!C��ڳ��..�bR_�0�3H|J�}�Ws����3�j��r���8�N��n��E��A��vwkqK��J�Pv ��2�t-_�Bo���H|m�y˹�]�I1������6t��k}2��T��[�-�,OC/C0����"�ɥ����ll�S	�=�y8��3�R�|�=UJ���=�7L@�)C��2������_8Ȇ[I(��$�z��dt�-j��.�\"!�1� �� !��s�sc;�/n�!�ս�@5��E�� �V�pL�S��H��t���N��jE�'B2' �v��c9�DK��y��Nn���9t�g���r	;�0�:�NdwN2��.޽2�z��I����$>,���AS˒��M�佬2%��W���oS2�]��
��0�)9,��[K[kM�>n8�Z�c�/�̱w�\c�x��b��7��d�:�W
{��D�11o������#m�m�
!�T�	5���Z.R�Bi�����S��D�x8�>��.0��U#�����}b�����$β�E�8/��4�A��ߥ�J��=�/lt�Z�F�%Hm����-3�W�}�����Ќ�ʝ
kK�#Ц>�����q���R^�Y�ޚ��'�s�Ɍ@KR/9�"T�=�����QK��r�����PY�����V(�q�f��?>����n��q�w0��Z�%)�b#-��t'cf	��������fH�>�!�Rg;1�?�]/z�AF£��:f���5K��Kfc�W�!�	�G�OL� ��J�{;v��
5Ϸ�z��x�ƅxV�&�r�c�%"����(5pL/64��]���!{���*��W1��[3:�:I�=�[e�,���hʐ�sH'}r�sSe�T+���HxQ[�f���9���Mc��h�͊����4���r�������L��#�Q���)�q��^A:[��N�i.�*>���A�ZYQav����O�ށ� ��$o�*��Z�2��.-cy���R��~�'ck�Ma��9L8lgܡM�ӈ.�W�n�#E�TE��I|P�#tP���v�����9�V��%;1>��o���Z�h�^�`X������{_����Qm@�ZAJ;}���!i��M*�/�T��2�p���m�][���)1��߹��y�?�4��*_��)
� ���
��8��@���.*�27Q��2Ԁ��ȓ��L��VVt�����a��M��>|ɇN��14�i|bq�~3��#K��`�j��ij�ɡ?S�%���oN#���;�+ݢ.
�*�)п�
����&��r�毠�cb�]7��M��QK��@�����96B��j!���i(�x����T��X��P�fC[�x=��N}Sal�~1�(=Y�����:�o��;؂���@�L�Rq.L�,����� ���7��b�:Λ�m��ӗ�#�~0SpC.������Y�B%��y�{�0����W��"^�U�uE+%��`^���<G(��5h�k�fry���� 8J����7��(@j������u�����94��
����X���ҡT�7d$k��T���PT6���;�����ܟ;���g$Ȱ��P�oj���'x�����P/m��fE��8�%�OI݊:��g��pL3N["bZ������6NO��Ȕ]2p�+��8��܁Ǯ�%���$0�0�)Z���Ű��U�'G�6���/� ��3� >�~�f�}7o�mz�h���fJ��b�=�/��{��
k1/��Q����=UF�V�zU��nӁ�	<��GF^,'^�z���aT�t%:;)�5%�����:=��6 �F���0���jlti �dVw�Xܣ�u����e��0O�����6�������C�LZ۲.V�~[�����U�O��926*9cE�L�jo���gd:V��*.EVf�[j��hP)�Ir��OC+ݹ��1��Qْ|�ν�3�Bs�oБZ��]��M�f�'�S�n����	���l߫.���!1���V7/��|!������s��s�ە�� /�.w�Uw2Ή��,T�έpͬ�#`��ͱ�=k���'�5�Y���g�$��Rp/sD�XV3LJ��ɴ͇ؒO%�gL�QU����JE�͗��qu�2��k� O�_йw���r�i����^�dWxG$� YjPP_0}��H1:Zro�lq�!sy��+R!� +�n�=�R����$��N�{�5&��K�X�����eT�f|m�Uc��Y�Y����O����j�ҫˌ�BH79Т}fݫ��Y'J�ˡ��"\ 1���ǚt:��I�L�L���_�MV@W9y��W���&�`���:g���+h/O�\�(~Y�d��S2ɜ�M�^���ꊏ��s��X�v�~�r�x˶>"�r��������0W&�|z`�וY��}����D�(a-�ؔӠ�<t} ��W�ܻ�ϭ�|��Ǫ���"F�3�weUb0�x�z�;�_dr-W���̀73�&:�r�)�w�k;����H3����r�\��~��Ҁ����-�FW�P�c�q��h+������Ku���q�����5��T `}Ǒ����Jzm(<%�����Y��_�m���X�پ��0�}�ٰ_��Y^Ɩ���N���x~I�ןgXamЙ�4���	n�v7�׎:����,C��p���:�
�����,5�YV���p���y�Qj�۔��حK���%~W�8�1OeL���[_�[�����;
֝�%%�[r~D>a���+�3��L�h�j"\ �.i�Fsyrz�0��C%�Y�3TGEǰ��o��t'�h��W����"��z��w�+�ӠT��&_1ti:gka����:���צj�q�o�]t!%��wF�y����ώ��]<i�1�YL�8]��)��Su�ς�F�La�����<sI�S}m���F�����Zx�K�$K��i��!�������qM���p/�K������Ĺt�h��{�d���E��V�j�����l��L��A��� �MX
�)��� 6��s��b���$k�1F��ǥ��+�Dw�كD#��A�i7ce[,d��X5�4��Eb�i6BS���0ਥ���ÍȿI;����EV�Q���_2x���k.Gj,�_n[�V��r�~2�B+�ũ���%�e����L��;Iʇ�,�~3E:Ze4fw�0�j�y�O�x�X3Ek��~ς�詒.�:c��������O!GJ�ǐr���@�埶+9")-�I��j���FC�Qg$��`Cz��Ih������O	
�~�۹�m�ӊ�m}��|h-DXy�D��͑�%~��#|{[uG�� �Ѓ	�F�O붸����6����#��~�ʍZ�ױ�Ǯ^���Eх[���ոۉ�C��V���.؅�	�i)Ƭ��ȚWOHj%����S���cСL��=�<��Yit:2�+��fE�6�e6��i7�pU�|����Y�	X\�bhg5��XA�M�����Pl:���Z�����{�]�}��XM/�)���]G���K���R^^�:�#��Qen<%���9o�\(3��Y��_b�h�� g�ħp����s<��h_V�+Ш�!�)�[�R�y�1��ޅ�39zE(H�� <����n#�׊8m8�e���7��іg[�����b:�3��³�Dl&C��[��\�̣���l�L�-�"�j�����ʄ���s�N����Y""����1tU4����_���MV��tj�(���#���oj�}������AK����hw�d7i�`H#������)�$����Kʬ˛�b����<)��X�i댷˵`�LG?�NS�$5`�W��N��1��*�G9�]�R��L�Li���&�Cr�wot�3�; ^��>�{I2_*�:״��_{#^�EVoa�U� �}�:*��7?�9�RzL;���=������!w�q�!nw�6j� �����A��qr뇼���@�ˢ9��������'d)��ܩ�q��я���i� ��װ��*����إ�?�c�	��FB�%8+��1$~�:��%�~�o\p퍧V�Ǽ��`Q�zՋ��=3���~.�#�I-ՠ�=]Y��4FL�贈#Z�iß)��V�L���5q��9D��@:Р��K.0�W���p8�Uߝt�3}r�$�|��̅T�+��o]���o�C^Q�-~�T�#CA���8���l��x�ȼ����4��-�<�����E��T?�!���y�����cL]�ӎ-�F��Lb�bʊ�ԩ%���%Rg���+�O>�.dd2���q�й�!d�2�U$|�G�+��������w���~ą�D��S#�e�Q�M����%FϘ2A�<AD1}�`A��7L�A& 2�����~6{��d�K�}f�/+�9Q���Q3�	�Vé� �}��2GE�*����f�.�Sj��L=;X��f��n����c��J�f&��`{`��}��31��#v��
tC�/�k���_ȉ��X��csף)����2/.6��5����瑊(J���w'2�<�����7�ўC�c7�̺@�޷U�QB>a���:�{աf��V �ǁ��<���n#�#/:w��)uM ��K�ōf�{cZ����������{��uמ1\tEv'�3?&�Ħ6媮r�Io��Q� g1)M��TV}m%�uQ���E��{�j���Σ�%�.����=��8�Aܮm�����
@��������c��9���-���?�K�u���6�[6�9+��	�����!H{`z /S���Q�^t��ھ|��mU�J7=���������M�h!9�ϛW��V��8,��J� +�g�"&؆��	J!,W����A�OcCp+Ǧ�V�ĝO��1��#$��i#e�͹�M�"J�����".�?ʙU-5[�(��ˊ�?�`�燈�If�8�9����j,V&Qoc�/�)��fnbO[\� tJ�*Sy�@����� t/�J�K�ϴ�:�]��}=%���u;����~aZ��|�+I�G����Z����rŎ\�X��1w'd�Q:غ�&��k�a*%"�����+7���ʼ�R_c�G��d�p�G�,���Х"G���)�GcK@��nkk��ѩwu�v�R��AG�.��+���ȸ₅�2Bؽ��q|�4��Os���%��l5c�E�n{Ӂ�#���d.o�/�Ǘ�{�YPՉI5�.�5>��#/��1M$�`#W��t:-;�mV�'i��,�!�DeA�¢9�8m����z�9�Z�E����ꆌ�p��FE��L�I�
�:�=�/Rb�atǌ�R�����aJ��-D�,�^�ǒ��
a�x/�o�L5���/W�ڸUSDZ�k�r�ǐM�r�������ɡ�K�_?�?�Rϵ��>x��Ɣ�K�,I�:��(��X{�R
D�R+���xO�2��M���e�
�����oYGEY��5�	��Z]+�{ǁ�)^?6['�>�l
[D�
��v�f�������o�q*h��`��=��y����V�>�<��<��N��r��Ql��{�8�������6��'�Gw���#�����	_ц*��ABW�e����-���-
g��	zj��CŹF"6�ī)ͬ�I�eqa�ى�ц
j��G�뼇�����A��cP7��O��\�F=79a�9M�$sQ6���϶�q,����G�}�2'�F+��}1c�/r>{� �e�N�� 6(�\hg���s�=��*�K���WQj�Lb�ͣ�I����@�����p�����4u��9�������lP [�yy�9P������.�+j�����P��Y�ȣ2��3��f+N�Ү~��T>�����}�Mj]�ց�6
/{0K�c�SpM�&D��Um��}q���/ڄ(���bot�玏��>��:��fyY���삙ȶ�|도�d�}�g�~���j��fY"Gc<3cV�1�z����#���.�P�5���IJ���f���+KWY~�H}B�a�Ms�E.o��L�p�}縤��M��cl\6�����v��0A6:A��P������H�����H��r11�:b�2�L~�� i�'�)��Z(�����}�(z:E��L���g7���n��2y��MM����Ch>�t�BZ#j��P����T�.co$N� �N���nU�;�z:eE���8�D[�X�~�g�\HN[�R~�۸T7����s7&(Y"3kn^ĭ�E]�;x-������{�Y<�����85��4�Y�*�Θ���7�B��I0���k=H�f��L���?�� UX/-
�T��܏���n�����o��F8��]���Eo2V�U���[��s�#߽݁�P��,�\���=��`��[�ǧ6b�� 8�"�����o�7Q�]��ӆ�z�����3s��W�.A�fok�(�9�\B ���
O�t$��[���ܹ�aO��阴�P�3���ρd�5��I��,6��A\�Wn�W�m�q2�� ��'��>nEWO����P��`8e�HW�'[X�a8>��e[��]��C��։�ծ������aq��a=����l�el��`�[$�|O�Ev�j���΄
C��t�1믺Ό������xڠ�(�����x�8⧴������Ÿ֪�r�H0Dn��
ܥ��7�!�*��6�2��P�8�Z�݊����&��!C����4|v05��ݫ��_*q^E�O��jC�_�ƜX��
���Ab_U�ɮ8Q8��+λ#/��zI9�T�QR!�n,�+q;�?o^/Í�^x'q*cә%i;@8��=�j[j�O+[���Y�`/t��E�og���#6���_����L�B�"��2�\�s�16�N�tn,�)<u�ff��»'� �j>�:E>oF�������<��^�m\��-��8f���l/i?Cd�R�� �b��0�٦gݘ��}_��a^3�F9f]�ٮwHa�YZ)M�8�;C�gx�y/��w�L x���#lG���R.��ePFH���T��
�x�����G��R�/k���&�e(�a���f"��'ɗs~;�$r��l��?���W>h��1D�Z#�4K�\Q|v�e��,�e��G�9!�;�6i���0������}]���Zs��|��/����0�i�ɒnyd�l�5����v¸ʔ���y+�8'Ā�Y*M�f�H� +ȋԣ��u�a;Y+����n
���[*�M�M\���x�K2_�}}UDn�v�)F:�AϾZPiA�T��7���Wg���-�2j�"҂+ɏ��՛Ӿ�e�i� �T��(2�"�곊 �C�Gw�����-A�\i$4
��r<��B��E�M�	]���1�a`�.m�сJU�������y�q������\{�r�ܗ�[�ygN�TxI����Q7�����)�q�ڮ���;��B�}7���o�2n�%mՈ(?�aM�O�Cp�)j��rZ���<����Q�.K��M��=>���*<����@����"��+y�<d�@����׀�=� �ܢ�uL�i`��@�N�=>���>��zeS��g;��>�Ӑvy.�둵`�y��|�.۰'J'�G9A�԰����0V���1���H���Z�8XuI���o��-;���$:P��^i4lM���?�cǡ]u�
dM'�
����L?V'`��[�4�*�:3��������B�S:?����c�O."� ��{�~_�H���QT{��yR��zR�yL0U$���l	d�l�K1_��>Q�<�N��;�0��~PM�!�|���C4�E(� �"�ȬkT�e��Qr��ށ�6�C+~���kD���*�W�\�z}l�F�t��m7;��73��4͓���;
y�����/�����%d��5d�Jj�5����Lz��z�,� ��[!S�P,��E�b�dS�ʳ���������+ӹ�b��K�w zԔ�d�X�V�"���-��>
v���
Ps���.��bZA��d��,E�Va�){VK2*Gh���rX��p�X��G�F����T�/�Y�a ���=��]pu�0���G
,�����0�A���s�C���,�L� "�Mdޘ\�t6���ĠcTo�R�����Y�$W��,�W��Yی�6��;���`��H8x��O��4\\sgp���7A�٨�<�9H�֮Ă��>D)^�3y����@y�B�)~�7�p�?3iM<�	N{'���P�̔晧����R���Ń���JU�O��Q��쮓�]���T�B�-f�~?�(��X��ìU�B<�C=1!�t���ٞ�9�dh�'׵�4�i�i�5�
��+�_uR�F��H������$	0Z�,�h!<^7B�i�Eõ*��w�Moqs�����L�2 �U���012
Vb�r���"Ԅ���Jb�Zm1�,k����6�����6�_��xd ����GgJG��h�0�=>6=�Oo�4�Y�Ӂ�#]uf~����l���^cԵ�8��� :p֊S����Β j��RL��M�Q���%{F3�2@�U��D�����_�fs½�	�|�1͵"�ݽ�qj�0�~�L�$�5�z�*&����`JP�<�����v�����4�̉��&ܘ*�ͩ��:ș����0˄�тr���S���&�Ň��ǃc�H�������#��������/�� '+7� $�fB�]x��+e�ta>[ �jݝ�&T�	%�4���#�š{p�ر-T��#i�]���A�U�dH����GS&�=����'���PNM�
lq��:���%bZ�TW�\%�|#w�72w0�U�l/���轀}tG��C�|Z)��hyx���̉unD/�$����s<����-����[Ǟ���.��lY=�oXK���e��;&Q)�9���M.���&�V�Z���!��DP�s&��k�G�H8�>�7V8�: )�Ԩ�$?��QP�o>����,� �:�@��8�*�n�>�R+�A���B�d9<�����vZ�ҿ�8��l�O�O���HnW�A��áN��˶�Ďs��L�lҟt!�
�����c�Qjd��㖕�m����D�yg$��-�-@f.ǘC���\��`��ղx;��T���+*5�D1���ݩ�6��(�Y:�hU�Й ��6i����G`���Џ �Μ��M	�̟S��Aԉ��]n�;do�k�����?Q~%͗vMĉ2���C���N�B�0���}�;`��1���ݜ�n��Z�v�!�F�)�#y*_�e�~׻S��@�I8x�P�D�T�'"�x��+
o�0H��ln��<���t�7!�1%�58[�r{&��)s�Ƕm�-삆�i��=�N�!���|��i�s�P#��s��%�\��2���d�TSO��T���a�:���
�B���7��;U����� s#�d9gu��aj�pML�:��+���!~1;�a���AzM�t���w�f̢�ԋ��C#�[)��G�}���5��?�?��Df��~'��D^w[���%�}l��(���F��u8�<�z�4��E�~R_�� ��#�י�&B%F�_,"����>��H�T�~5�4ы��k��(���-�x�U�b�g�YPf��#�Gȇ"�h`��:�S[,	7���,�� 㔢!�����9W$��s??�u:��������چZk?�ؚ�`�6g�0�[�aʎ&K��>�徴(�Ŀ�x�����}�M�)�!�"|���=Q'���'�Y��0�W��.7U�U�/p?JK:�7�4��ĩ�@$��L=r��~�2� q�����m�1�s0˳b!o�5��:��8�*�R\��F*�)%i2�r��~�ƪ*��}0�-�U��Ji
YR�i�ݴ%���)J�_�; ���}n��������O�=��A'_b"?�E�b#3
Zu��Y�X�V&K�53��v-��,�1���V�I �N�"d�1��s���N����<*�F<� �9�qҀTL�@*�7�����z@{�;��'���s��V�Nܼ9x�����Z]L�KD���6��W�f�k�Fc@��x1*���\��~j}!O[z)@@W��O���<h|���ɊK�.Cft��U��Α�v��_�~}[�X�z��k�=B�cŶ��օh-s��Ծw�h�^�bN7!�4��`��F��CT�["����'3�)=R3u�J����e�ό�̷�qǛ��'�I�}�]���8/oL�T��d����fD��DƦ�dt���ǐ�x[+����MO6�-�8�֪���>��᷇w�ٗY�q��Y�=R3P7�e��e���(�̫�*���y�<m��=���㽾����od6}������U��+���"K���xh��nw�K@x���x(0<s�ԦvY��rI��]-]�a56W�u�?��'/�8���Y6P��W�UC"��e�g��	J��/�fw{�`�p�'�%O��4*�NHS���hP@M�O=5����W2n�뇤-��`MB���6�ڼ�a�}��UD��0l�͆����Ç�p�j_��V��0g!��֋�����;�;9wzYp�\���0��/�O癓 �/��,|�jR1�,��z�|�8��2[���N"30���|B�3��j�D�j��l��:>��D��`UHX���/�Ĕ�4�G]tDIj��y�<�k�6��&8!��Z�����h��� ��4�����3˳-�3� Usi�Y<Q���V�ʳ	b�� � �����x�hyQ���.3]���!Ur�� �q��ǔT��� �LE��X�sX�n���n8�S:K�t�b��~�VD�-�#A��ő���n� [>�*o�\�ۥ��GK���E0�;�Jϔ�qp�C��좃#ЫK�ȃWE�TU�����U�V�E���z)�t�Av���F@�p^ �G6|"�ۀ�'���!ɸi0�s@t//'[fm.� s�H�]O�Ϛs�Txݽ�B0}$ O��I�0�����bd�.�rjW�v>ᨯ�0fH���fB��f���=���ڀ���Z��}~�Ӹ7����,�8� 3"�A�b!i��!�dx�߹�~o4����`�͡�68i10F�d�r��yE
�n3��D�H��=�r6�wo%������οvR��N��8*vY|/!�Qc�e��eu�� ��tu�M�f��&]_�A���s��}��?�vvX�������)L��xAE��y����S�H���ī�M�tzU����	T�n�����DI��ȸLѯ��;R(#��*Yz,,�wr2v���:�w:������d3`H������D�cX�S�j������iޠ�Ç��'C�A@�a�%����C�Yj�w=���BB���G��մ�\���uO`o��daz��c����� ��dnE�`��0�A���ye�&%(: �\�OK���ލ̙{m~�$vKS�e� :��x5"�
����Oh��N�����9$9���5k��?�(�+T+��XK�ɝ�3a1��`/]���R�W��tn�I��c܂�X�I�i9�u���2���x��<f�����?M�t���};��W���;Ҿ*R��a������,��A痛J�V|�Ɇ���f2�����W�u��h)�r�!��5�~�Y�+�!�K�I�u�����%F��S#�L��̏�[�0p��z;H�v7��c~�P��UI&���M\Ѥ��^v%ǟZ��n��%��a=�L�����G��uP��6����Z�uz���H�������ſd5:~f��X@����nM|$�.��R��eִ��T�8�!l��7u�<*�
��®�M�YX��2���A�}�v0y�E8��6a�v��"��`ƍ)x���p����a�P�D[lM`��QD[���� �㷏p�4L�Ħ]�U2X3��Ju��R���H�`���ל.���B���x�T��ǡ&�Y��gI�uY(4��l�s/�r�Z��v��}&�5�%���s�z���ㅔ��uI�]� zݳ<z��ݸ���)��xc��ń}�%#ϰ���h���BJ^Y�X!��(8�
�%Z&��{��.nR��w$/iw�:�r�z���df�v������(��-�o"𹗛���W�yP�j�&�jt�z�O�q�~���g'��"졡� guK�tîC�}�u�ݕ�5h�`�Z�T�Vvy���ܝ�v�����Qƀ2�z���(�,.G��]X8��혎k�D`mBXa�jq��|59��Ԉz-�*��)c{{}]�_K���=�e�������˦���GxE���ѷ��8f�)=�M����r��u�g��AI�	x�����q�?.{��'�9���K�/˸;=���Ǘ*���u.#��=��[r)5���+`-r$Z�?<[��	g�"�+��GyaÙ�b3��ho��V�t�z�����w�m_�������@ՠ�
�wG����:��������-4�c{�w=.[�U3���M�e,��6���(���+,�]����Q�p^�&h0�H'�,�X�����"]��z_-�0��&$k$Z�P�Eu��F��n����Ds��E<+@��S�3�[*N���[BX}��5�~��kk�ą��׹���V&��蝴�>v�8����BMqB\+���|zD�F����B�!\@=��ۊ���y,G$�vE�4�Z�Å��i#ب�^�`��!ƌ�a��nSp<���x kr����|J"R�?�n��� by0�q�L��}@~䩹�f0�S�������`�z0nZ��k��.�\�%07s��$�z/�Y���븁f�E�WU�B wқ^��)���Z����o�A���i�� @ˡ�0@ c,���۪�҃��,$�����m\�=���x+�=�Y�P݉�ڶ���7T"�h�$�@�55��Ec$�0��)E�Z=J�j�$�'�[�������W�e.8;��-|�#CY���,7�O�E4<x���0^���F:��\L�?��Vp�	%1N�
�(rN��qu�������pk�!��T�	�D�;=G���S���\*+���a�|���[Of�;�~��Hj�8G�RL9�����U��g
R;f�����*�Y0�P��'�E~���إ`o��k�2D���#���E��d�2����
;��TGN伖C����Z�I�p�߷u�3Y�+��)~E����xw��Wb�0���8�84����N��~�x!g�9�X�Wύ#�A���<1���~yos� ���\M����y������7� �M��ƹW�a9#�v:&�<�8�&d��%��xؕg�o������[U�r* ���[t�f�\7�ā��nN���P�oS��i$$���`���N���W#[=���	Q3��Ludn��o��䷭���3���z0�:H<~/���b��ΰf��Pث�5]�?��S�H�й�n�*�|�� �����2������)���)��ڨ$�X�w��x���R���D���7�]�$�k@�N��ʧ�&��iZ�Q�Ss14��y0���N>A�5=�h��h�#I�F*!�I������!K��:�+, �D$�C%E=�y �͘���n,�"�G�4�Q�/���'$,��Ǳ��Sے)��e.�PJ�N��k�j8M�U�1{����=Άo���+K��K�Qwf�}o�n���$�v8Ҝ�/�㉅f����� �&��a�S
'!�m;����5M_尛��P��d/&�z
#���D���Ĺ��x0.�HМ��ʼr�rd4q��|w�[��>�R5s"؍���X�~����S4��f<pj�����5��]N�N�,&|Z�ݒ�
� �����u"��Ϻ(=c}RW^L_=ށ�~b񔑍C{��x��=�pp�H|o���qvB���y�Ƿ��1��,R��	u��x_S��ݿzh˖߄B�["Z���G&�m���.��=жǏj
0I:�f��Wc=x�/��$�f�mw1���*�:��J>0m[i�H�8S�N�yC ���vԅ���eY��	O�@$C�+>Re�o
��c��:���R��B+�»~'�%Ẅ�s�Q�"�N�4�A<����m�B��5@����N�����!D�t%��>u����V���v�e��J:���� ��c�0�(⌞�7��*v����
6�ڐ�Oԩ�n�p=�Q�I���4�B��>'�:P����ԟ��Ͻ]���Ye���Փ8\�Ph�j�|b4j7ώٳ��d���� i���JW��|
)�uf>�a��#��1g{��[X����!�Dq�<��H�h�*
g$�k8��B ��x�Lߚ�� �����-�e�I'S0��\uG�L2#��t�x��BAcP����� �լ��z����-K���0;ܮ��hi��C�~�����Vgj�4(�A!�2M��`.��,�@�)yr@Z�v~��T����TP��qko؁�5�i�6��	=-��=�.)k+v�b���M}�4}D��i�D<FD#���<�O����\6������MB�ǫ�����_�~��ýMٶ�WX��O��u{3�R�+���ѓ�F} g݄�����D�>&m�M�8�B0�.���8�����v��h�4)�� �!Ggzޟ�r��P�����e�@xx����dq�g��W�@s�q&Ćc�Xg``�b%܅���"mޥ���>��˘��t��B�R���[�-�����!��s�ϛ�j~i6�6��Wx�ͦ��V���$��ŊT�;~����Q���a��^3�j�"6-�i��KMr���FB���W-���p�l5͢��DJc�o�x)�GV�`	�79����7�y�"���2�� =Z����(x�.�&I�=B�_��>�P'b�@�����g�J���@�SƂ�����H���Eo��$
������%�؜������?D�\�� DM�����'yK�CW���,�a���yS�e�I�+]|C���BR��@�d�y�����`4J?����B6�GS�*c��D-Q�^6`���$��J���_bur��?���[:�tz�?�k{�٠ț�vrm�C^����t��6�����e�.<J{�p ܽ
�z����/D��#H�y� \pۯ�D)��Tu@=�׺9���ō�XUoM�Q����H�}"����qR��,��[�_O�
���R��17�λ?������w*�Y�_A�~�PTd�B;� Ȗ*����%���؏ֆ�k*(�P��m��~����4Z�Ӝo�,�VWoI��M�nzLI�	2�+C0O $�؎�Z~�n�P�[E�=�r�\~B��g���е��v�K�-V7�'��-HB�U�E�т|h$����7жk�c����@��wZ�����R.Q�	C4���E$�d�+��}�<W��g�E@z�"�l8_�"%��&fs���}4�`ƅ�LA�$/� "�Ձ�r0���Pof�t3��IO��u�˰�[��z���U��"�ֹ竲x�Rp��G� ���K��E0��t�j �bq�L�z��E~�B���΢�*�k�}b����T�8&|��?5u��/!�),���� ū���M�f��OCB��ǡ;�4��ݧ�����K'~'~F *=6�[-A��xF���W��� �ֶą?�^%#�b��/��!&�g���܆n���A��$|���k;�I��&��k�v).Y؀��+�Ys��Ejt%h���i�B�]W���_0�N�(��y1Z�"����������QBn��'�x��6����!��X��6ՠ�{��-=��H�M1"��S��gv�>WAy�x��땠�>�ND��y���T��jF�%�t����:�+؇�G��B��!$z��Y-hI<T5�IK�9޴z�@�+������Ϙ
,��M�j����N���0W�,Gh/KYu�f�M�~������{����,�Bh��B�����I�Pe26���o�߬��XG�TmG�Wkh�F�Ab����ظ���fB⬢b'�g�5.�D� ��0> '��I&��0\�tk��Y�hg��O��^�(����6���IE�$ȓ;V�f�Q~���3�e��|�Ã�[f��#NR�nіb��˥�X�VI̾C����=����r��G6�Rhf3�>�z.W��!v@�J�P[�>vh@�g3������*�+Lc���m�e-�1�Gi���쀋O����h�"L��Wu��F�O��DT$�]�Y/z�ȷ�.��QI�D��?d%�h'�{�{a�T��㘹u�����0 ��X͆A�al�}�%�L�>�aP�x�����+Z�w�|�K,ԛ��F+8���4P�3Ol9�ϱu֒��e��y$������",Z�~m�\&����PJ��w`w�"�r5��4{q���#9��s��$˱�����n���`��VJ�h:]�z�"��;���0͟d&(�h�aa7��=Ȣ�{���l�����t�QǪz���诨pO�(��U~�����j�מa-YX�g���2"��02�1�������:�����:��w@�:DS ���Хr�{©C)fÅ��q\7�5�[��Ц\x<(q�~��B�>I��k�d	�<���6	Kx�-��SzoOQ�.��I��aș���r-ȁY�s	�Fy�w$\@vz-b�2����ξH���]�uTt)~��.]/�ԇ���l�}�&�����:�8����X���R�����&��?2�$R�۟T�X�P��lJvl���/�OĄX�s�Y���1��=5A���!ǋ/�>>���#�DP��j��ya:�F���[Փ��?�/�a��L �S!�?)�ۼQΪ�3Xnbt�a�*�G&�-��sv��n�)�ݞ22�П�*�9��ׁ븦����w@ J�4��!�r�����/f������u����m�o߂jmD�v�h^Y�(����l�#ݜ�w>/h��WK��mt0�/&V�:K�xs�o�8W/kֶE�	�*?#��s�%�������D��Z�P�E��Rs�j����9�qw&�^G4)�����sC�	G���ߒPQ�X�f�alH�k��B��#A_��o~�QHMX!2�Z�^��(�>���:~�\Ȏހ��� *|c��%��-�耶x�k��U���w�x�+���s�_�/*�f��Yϗ`WR��4ۓR�G澺�h�������Ĵ)&�v�8R�Ӫ�Q��%ͺl����6����q!;yHj��)����>�q���"R@�d �$�۲X����y�6��y�|J!����}���ዣ4��3���0E%vP�6�v�D�v��w �֧�"'�gb��j��nM�#;�o�� -����;�$�u��!��1o��p��O�t�\�n&�ʲ,�ٵ����>O4�@�')���&�q]%������lTP=�>���v���`���5�\i�}�$�q��4��Nj��<[+;�P~1}��dRS���t�\�^R�>�ۄF^�����"\T�J�g#W�h�4=6�W8��$c�S&���bo3��X)���`��+f{�uGKآ����� ���N��݅�oZGlAM|1%�T(ͷ�l���K"T�hs2暹�uٱ����;��(�8g1��JQ[:��\�W��δ�'Q�0\ƾ������
����#칢�]�w��N^�pP�?K�����u�w�� ��}����`	��2�������Ξ�k 	N�̻���:���m��t�]<D�p�V E`��Pp��_�&��&ƨ�����"�h�MC�����ww�����{��s ������s�uU����W.�h�&�P�F��5�ϕP�=6z��z, �mm]i��b9�c�,��i�Z��@�e-�G4}%�-��K,�����(��N�h�X ����)�%G���NڨNUQ�ۄܬ]��7���%���?���O���q���$_��q�0�Uw�Ni:$&�.���㓣&j�C�'����s��Q�7�T����;��
���4�N�B�WpE��� 괩�3���KV�R�a=���m��:����󱜙/Ï�p�j�}--?�=Wr�t�y|�s@*Ꮫ��mK���=d �.z�f��U��$#��@�B���ьRp._�l��Al���z�`h�+]�Ρ�!i�6�[0�B��H>��H�ִܠ���'��dAx�X����&�מ��\��S�d�E{덳�62��t�#��U�B�����B3K3C�M���rFQK�H.#m��EV��<���$a>UI�+�c8��ЯUCEè`�u�L�<x�?�ϭ<���6��k�t���iB�o J�7�ש�L�1�)s܁��iV��@���2�r����|4�S�0�GB��曺��=���kL�pT�s}��hv���C��B��8�''��? �3�L���ns����:;㿧N�yݐ���]ŋ�릑��/�l�)��;�	�6�b�"QL���Ka0�~P?Z�h��q��T;b��7�)Q�ok(�8Y
:�8�	*�3+e����K������u0�
V/.��M�z�]��⤎+���������].�H(g���[av��8��萐�E��)��FMN�A�`���ά_����pO�B� �õ�Sķ�d2B�smS%̜���s��qd�b"C�!�=`��V��H+���b��=���3n��U��K�X��`� 0�zznY�v�6�q�v_���=_B�H�R ��9=�{hO�Uc�Iub��� �Q ���R�욃e�rǄ�[���
;CH���o�fK�e���ԛ��&$�'y�s�N���:9���l��}�ի;C4|�:����
��?)��Ma�ѹ3�]��߿�D�r+������d���;Z�(�^!{T�"����[�2+�T[�8��w���o�:iե��
�[����z73���)|k��.��ׁ��H�׵�q�]*we�Cl�ɡڢ�R���ڜj$���X�Ӹ���d�	_�D1�6��tx�f�ʦ'Y6`0�8�l�.�� d����+��0$��b�]	�^ ro�y:8����ǻ�� ��=tĩMhd�CP��OIQ�֞`!�a��f�f�6��+�q�����L�վS˩&�+�3����Z��' oi ƕ4_ז�I���aqE�bfS槌v��I�P��p{��4�pz�%,@��2��4�>|ūR�Hv2�!�3*��1��6� ��^�LI����:��
��:a��8�{�J�X�'�,0�8�o��.�2��
���?�=���\3�W���:ˎ��k��W>7�vUo�vG�J������ԅ��Ж�*��vZ���˳�чS��aj��^�)4�P'��?]�+�̱yc�0|0�*����+E�/tv�w�r��E 3.������rI�����4�z�_c1)�a�ٟ^�y���M�D�Ŷh�*8�y�}rh����R�-tN��	�{�:g@�z��S�ʾ�]+��FPL������*z�Z�� �ŨQe�IF�����D��"�U�5M��N�.�PA^��:����T�&�3����j��o>Sav�4���D�=X�0���޳s�W��1KA�o��Y�K��Hy�_i3�k�zI�R\�p���/{7�B36�j6�9k���{���e��j3N�g����xnN����m�ϓXM�6{ަ�0��lt�	�t�z�b ��,�Q#y�ɨ��I��aw�m��.=��@�R�t���L�fM�u�Z�����J��ᗁ�uD����J��"�2Nh-�'el^ݟ&�nߺ�����1�-���}E��Jl�ys�G^ˍ��$P?Sl�}��>�9\J�Ǹ�W��|���g�f�X@���C<2^Ŗ4�&���~7I%�rb=����{��Ow NT�eا��<��껦�r�Qm�/2�r����%����[�ϭ��
��+f���W^>=��5�V:�k��!�s��σ��Җ�����u
eńl��`z�u�'�vC�9i�bJ���>F(��̌�ao�]���hA���ߣƭz�
^��{,�I)����[�k7Ş���bf�����́�}��]�;,drvdz欖�'Ba9�;�Y��F�Mr�X��ߥ\��.�=�M�i����Ȳe:����Rf��1�&���u�Ʒ^������1)� �՘��fF�t?�O�cڎnF7���\����a�$�4_�]�<���L!R`��C�1�p�C6�p�zD����W�#����AτD� l�<�����ɗ����uc�m��
��ǵ�8�����90��c���ʈ�U�-�V�y���-SPcL}�-����:Np��$�Tc���a5��T��D��� 4pJ��\[���1a���t�`[E=��+��F����AޞLT@����A���[t)NuN] �>\��#_I��T�Ӝ��\ȭD��&�!VL �ԦX�O���_~c�u��/�]8?�����Tut�Q�*����9{s��;�j�"�z3<ށ�2�A��BWst�n.��(~8��k Ί�s��I,���\��{i��[���ث�D�IM�⡇�1w$|�/}H����Kĭ~X��@� �CI�%���7�-OLT|�*4�:�U�?�r�u^��|u�# ��K�U\�t�䎯��j���ί*��m.���U"���-)¤�-�jVD��Gw��@'�2D{D��c��*�6wC���/إ�:'k8l/�lr���}'5ۋl�[��(�u��rՓ{S��N�ekNh:��uf�������:CP�4M�s$�{s�7HqY�֠�ʐ)T�֞�X��¿�N�$a�,?�����,���cH��y2�Ymt��m��- R�	��yPC�]���&�φv0��h��SC$r����[j?��]x{g�;h3G>�-��1��|��q��5+/Һ�,/���b�7,��RC� �����tzfp���7-1��"��g��qv������;i���Rw�Q{�dSڵ���"m���6��n36�˾R���7�i^�2BR�R,��h��4���9C�>Pe�OV����/!�
T?�VJ6/O{�b��C���C
R�X�O�J1���]���u��� ?�5N\>��D�*5�̈́q��3�I���hz?���7�L�ح��F\yӡB�K%)[0�h����k�3(C�>&�����2�p�-6\M<�[�� P#@Ň?����<�YN4*Gj]BR@�[���x��#�{ �)�0��i�	�WqF|}��s�5�Y����>ߎp%m2=�4����P.�|Mr�`s�	!�ƌ�@l&��z4�.C�	�e����0�C҆R}�D������b�����T��308݅�9v4�t��A��?@�2	/�iwܳ������G�TiS����Z�9��v��IZ瞪��G��C^}�o�6+�U?D֋-��x����wP�E� w�x���7��.o� H�����b"a�e >e6�W8Of9�|��HbI�Þ��ȍ_lc��[�49*�fjJ��Tkvp�q�@�h��s�iҁd����9��r��o���>G ! Rwo�y�7��s�@� 0����ȗ�Q������8���C�S��G�5Ԙ�`|�h��I:v{3@���p�l���j���J�(�����E�ZD��Qi�ʛ�ĩ��%p��#�-���(�MUMД	�[��������+�~�'�_���B�k������è��>�e[	N"_�ECY��&�s�F:h9<�m0�6Ց^���w��
@.�h}�#���G�P�صb��H�%�F��t��jK�gC���KZ6�-�j����6�����h	�1ST����L�F��K�*q��6b��uwk9��&o=�l��}U��k�1)���;D?�#4�5=�aM��x��� (��X��Xy,�{�l��B'[W���ES�?^	1&�!���R�B_*	���c�S��
WC��BO ����[�>s�%����w	���^S�
��%���ka��]r �&Qb��j�ڬ�BO����J+.���&3�������\)EJW�ȗ�����9ζ<����җ?lH��^(�����������q{<[��3�~���@��f�^dR�Ju�\md��]35��S���>�9�)-�R��c#p�4�~ 
}h��/�1}����|k�v�
\]:���q*��f����<@��r3w�6z�渚��?���L����4
.��3T��tX�2ڞ�����D����+�-m�i{6�1�4@�|����da����'���?�;��L^T��xs8�Ia�)D�:d���tx軠���#n�d�JvY8\-�6�������Lq�<�.�;\>"rVI�� ��{�])��|���ӖaO�y�r�mi����H[�e��� ֕����z�����:�\�dҶ����^5`[�L�[��?/D�ύK��~��`²=�.�S���Άk�L|���+�z� ��U|���K�4��A+�J9u�Ĩ-E��g�ȩ2��'��wh��ZF�l7��dsۀ�!���_��z��#A��F�fMg�Z+���9���7�%�g~��e
����K�xǶ���-/�%�S*kR�q
��%՟���B�Cy"Z����YU�a/Ք�����~���f����L��'$�"��ٔ��BuG!�����n�GPe{ ������W#�fO���P>�z��}�"\�H���6�����A�.�~�u$8\�m��ï�T�M4����3n3��H���.��+�2}�4j<:Փ������yIo���ݔz1��,N���~B�$�	[�h��{�B��)*+���r��k�D�=�iH��;uF
�rӚ�yB5v��z�Z�9hC��qu��%E	�|��w�{FR����=�?<kǔ��LD^F����ލ�0}�L{�B�k��Ef���T<���2sO��7��@��x��R<���NDHG6u�^��;�}�
ȉQ	G:)��&�&�p����P
��� ��Y;�:�O�
���j��ѠV��lF� &P������J�����6�@b�AB�1*�[�%�|%_47 jw��
dn~���(:�G1� ��Tt�xL�l<+���~"'�����Vָ^�!�]u����%��u6���(��v���Z��O~6`�-K�	��ù�{݃K={���^V��-�v�]�s#�T�c�<�U� �L@�4�-@��zO��kZ�3�D�5eE���Z��
��z>d^�"��Y�1'��d��S7u�U����%m;	.hf����M�0��dQ�$�ehz`��~!I���M�9\�J�;dH�-�Ȇʬ�s�YԈ����ɩh0R�M(���p�ieJ��� �%k�2�
J��!n]�����@����5oO'�)��;Yx2䅳�$�,�d���[�~�,2��ɗ咼�q�;�+�������h^Q��x`�B)��!��C�~W�V+���M������ ��@��E�e�mHbǏh������l�������B�����{�&Xg.�5�j�N5�]�<���mA&:�8ӟ��MǙ�]B�7�7e��^ߕ?�vH����ю���~�`�R0~b�Q`�� �������-ջ<_)���U9�l-�.ҶP�j}���ǈ�\ʀ�8�Q�I�l��tɘ�j�!����qL��(�+�j!אb9����y���J3�&�ƍ��P0�S��z8FÔd��;.�h��i��X]4+��\�<kTfU�XS6 �1Bm<���e��d����\��	N9����4�l��o�����!����u�O�fDl�D����:��F�$L�$�Y�H�L���Xg��H3�j�R�eX"/�k�~.�+����=��s:i�3q1;�O�X<%`V����qc�~�>p�m��t.��H�L7hШ ̸���ۡG�����B��i�}Ђb$ޏ�H'0��jH~*��0M�a�^@U�婞VHk|*X��D%���v��U��޷�}��湝e�0N"���3柆��E�u���Ǵ��o*�S`�ܗ/�L���$c^D�db��vb�[J~}:fwCM�^0�M������!5J�|�~���0(��>�������&��#{~��v�1mE�Z��,˰��x���e�+_�ֺ�ʅ<;NW��mH�s�+^CM���6AI�)x~Q��k�d+�B��V��J�M��������3/5~��v'��પ�`m���H饩���m4e�`�!^{_ͫ%}�ɽ�\����E��L��=;/Jl[Q8�����VrM�z<�R��s˿0�n��҂�*Z������ߚC��T�pc�i�ƃ�����~�T[^ڵ��f�'Q�?V��Iೈ�5D1Z�BL��%�t.# �@̡Z�u�z&��;~�0Jnb�����LBK����ٳq��_?s�Dl,i\�#��\0Q�&��'�r�'��Ŭ��/tO�0�v%��%� t�'�߄�tc~�]�0���ا��D�=�ƴ-Q���R�Uځ1y�1��j0܄�x+TΊ.(��zH��"2��jtl:61b�`���k'p���y��P�%���@������G>�-+=�0�&+�*�C�#�q�
H��_	�f��
���Y�2���nw�>�Y���Jv#^�	n]<\Wz!ܘ�W$OI�жq�.��U`��Y|,"c�61�&\�����h.%m��Kf2��|Ms���KTi5��3!����6$g�ƎῇL a��0s(\_}���ƽ��6�R8�RʳQ�ۀ�r��
�@�ê�y 1��O�	O�g�+�t%z���"����C-�
 X=up�]��9����8�ꖘC�ݼ�Ƅ�n�c͂��W:��{�N��@�B�d�������<��tQmrV��Ʉ'+UY��Vi-F�a�wkQY�D��7H{�s�����*��`t��^��` ٳ-лF7�Oi���u����#/�}�_���o���.)A쩑�B�g@�o�.UQ n`y�9}w#DV=��� ~Ϟ��d�nn�;۵��e��%�7nO��$
3�%/s��յ�$��e�A��b��,�[s�q7C없 �)����;�$Ő2�Z�k3�0��*P�E�M[�� ���E)c����a��ukV�r"�д�C���s?�[�Aֆ46����%��\���E"�,;�nu����#�ۄW@h����^0M�=<AP�W$*��s�ve��6Uo�vF{�BV����д�hK�y��ud���?�N�Ũ:�2�%�~�i�ļ����	!�,�-��ڻUxP䑆P
J��ѳ��� ��a���s�W�i�-K	��	Jyy�b�bdʶ"�#/Ĭq��ϋ=b/>����61��#����D=IA�ErB`������P|�n��쀴��dE��t�A`\�9V�˽)Ψ8�0�wM�A����XFˏ��ݘ�T�U���%z�U�h����^�����3ݿ�^����>[�!���O����Yۯ�P���m�"�������-Mq���5��C������ �4�u�3��R��1;=���P������f��(���کxdq��#}68��Wټ��Ӛ#p���9�X��6:p�o����3о�TƁZD�GFr �}	���&r�g	���B���VpM;�H�΢kVg��F��Kq4��?~�h/Y�,CE�0����Ynv��"|[��
�8��LӀ�S��]��ېf�^�}�n�{�T���%BE��&���r6|�݈�=��}�u��&�ܰz&������o�f5z���q�L��s��pw����k�7?��1�ŁM&M�����)��UY��/JW78�[�/�7�h��O	�sI�9��T��	)^��~ u��OQ������?���1*�d6��הP�5O����ƷC�9�7�;�O���<5�cO��ei'c�~�[;+���\[nͳ^�>6��-$%ڷ@_��a���ipӚ���=#�C�_��A��\�?��{����S�[%�� �B��ڛJ��봯+Kc��E�!��mV�H=�սל�Я��]��}�֬�~���B �o��Sgi�����c���"��*z1��1tz�3����4�l�Q����6�#2��۫T�: y���Dgю����Hr� �UJu#>�����LT�1:A>�^g�� ���v{rȡ�÷֬��h�Ia��(fٍ�Z3r�VC�k���l-���� ]���KV0s�:}Vn;z��FnOU�z�kْ|���)�q��EJ�ŗf�"ZR�(u�?e��}e��f�7�]2BFخ�;CCm%�\�F��}��z�o����:�{��_5K�^��^�>߷QNɽ��#BONSA]���Ðd��o�����:�H��̀�M!/�Ð�e�������P0��Ԝ�d��j�s�b�?ېq1����,�-���q�`ڐ�j�T�8R(���$���K��Х���-�r��˓��@���S��
�s�*N��qT4p��رS�-[��b��2� Y��W�Qa�8:���?�ҧ�/v�"koe�rfV��|;Z�4�� �m}�j���$�ɑal�帹��`[���dn��^"��C|ʳ�5i� ��]:͚�
xw�
՘��;^�h<�#7��|��b��_��_�W��rX�<�^uJ_Aw��Q�;@-T�E󌗭9����0��\�Hǰ�ڏ�����SW�Q���z�-�C��}����څ���zKN~���W9S��wZ�q���#�*j�"�]͎E�t�����Z>���s&����s��W���4(Ղ�΃]��,����|�� +	�,Ӷ�n�7:pjy�%l@4���3�Ʀr ��㙔�p�����H����=e��'�qdM	Y:�Z�Q;���&��� ��˞�.�7��mjѯ+|����٣�I��d���bV�Ě:ջf�X�SE��^;��D*,���BO�V��+�5�\��
�=�D���A�o�_"�>Of1��h�q�xӉ���L &m���?�Bb�,���p@X��hד'j	�JZ�@��&o?�P���Y��C����u2��(�F����	@��VD@0��C�ԯK�8!*1=�\���'��ׂV���o5L#�o�g�.��1u��3h.��F0^-ﯬ=K���{�U4l�����AL�K���Ƣ
l��4p���,F;7Ģ����x���U�C��������:����.�`B�/$�HJg��ȵ2S������AՐgK�N�Ǩ]�&��
�-hqܪq���ǉG�ښ�I�k���^�dWD���5�p�\c�0b�D	�mpf��Ѯ��\�iIĽt��"rO8�X��w<vnsJ��[�/�,E�Jʫ[�0���\͔D���w�z����L��L��� �h��:�K���g`Fś�������c6�N0�������؉����`��H�rk4���KU����*��T� ��b� �ʽ��x)Ya��u�y�X���/A�B��t?�������29.Q7�԰ć�/�Y;���G帷�#r�\��������(�?��m�>���	-��z�z+���Aη�0\BU��.ӏG^�����*^���v���b�DR�u�X��c�Ld=�'���#����4
�v1	0�|u�F
Ĝ�0F�p�����h�������0f+��ak�ڮ�iEt��E�,��f��JInpQsd��(1�^�!M�I�6���O����rLHXE|H{[��H��`�ϟ ���E�ZE���ݩ�:L{M%��i}����b���P�b�PR�<jo�5̹׈D���l�jA^j�e���n
�FY�5fَ��},��s�T�+�nw��������i0�H�����k���`���9T��ttp�+��fOx���(^'���B�^��l
>hCT��4<�dl��ω��5Z�?Pݒ
��Qb���W���x��M�v��3PaƓZ�9SUP-nq�.��_3�����4�j$�J擇�1E6}S���H\���Њ�������Vmߡy�ˑ��`芮�N�b�0)J�F���܃[Νc>��I�]��5�g�D�7x����B��/�i����1쬞������e���&@m��]��AY.�5犘t-��7�ׅB2S��[/��T�d�1�|�-�NLS���|��~GĀe�f(��)#���}�@�F���|_FU�%�SR��r�'a/�딁g�rör�� r�+G���G�ޖ�u��p�E��q��0ip���ţbfPD��q�y\x0�QWď,0�/�/�%l�)̂�FwR9��^fY-�s#���[�~�ʏl���2�̎a��3�job�b�M\�tt�����ܮ7�ᩇ���_\��V��9!s$=.ă>����p'�6t1��;*L@A���N'z�-�C��{#@��My�`+6�������r���h<a�j�,	7�R!y�����t�S�|��$��zA�nr��1m�����Nv��F L�__��|�L�<��
��6���d��Q,3D5���Q��I�з��5�����|�������f@䎂��e㴒�c��12�k��U~L&m����Bv X��==���u�(a���ٿ₧=�y��U�����Y,�����%��C���L��I`�&��V�{u��k�5�jxsM��48����6
�W��ؽc�٪}�}�N�s^Y܀�m^M��8�V���|a�h�7��\�PE
m���#,�Z��'�ΥB��D��|ވ��H)�-�\i |�U&����=�k��������U����Fp�eM�x"^�0k�1��{�Xצ�)��߫W�l�f~��|s&�*��5����G���B�`�(�S�D%V�/���xHT��1nƆ	ʋOo�f	v����y��e
.���~4٣I"�\���5�_��'ݺ>q��r��ٵw�c42��K:��Q���>]o�˜�h�1��rC��Y��[�ߓ����ܨ� `w6��l��PTr�v�yV?��D݅�!��nh���q�TM��C~+��(;��vT}Ȃџg�^�2��J��)��k�*f�/z��%_>#�!���.k��B��S���?L�)�C��B!5Eڭ���brs��kA�U��(N�� ��j�`�O�+�ߞ<n�k�'��T̴-m�B)��$�I�,�1Ey��B�n.��2���O�>���묙!�Ch�絑]���̟%��\�O���t^��n�ֶ��k�xyh�����P�'�߻b��0~0���/�hl�����q�$f��4�ج�h�H-F�QN��yc��d��H�P<��2ABM ��$��~�0T�/���5ES��V���3�!�0V�b ��������ׄ�>ei¡�-��߈8, �� �>2]���A��	�����oï�P�Iek'|A�/Bb��2E��V�S �%��]�B'ڵ��r�a�����iJ=ų�B?�e����D��[S/M��W�$�O���/���[��{p���Ⱥ�%�mԃ��ϑ��y�s�T1��Y��L�:��g���j���V�'xg��Y`��H"�Y�o1B��� ��CX��4���F�l;�T��e� �3�a�&{��z`?,uF��l!^�ŝ�F@9��P�TR�Gچ�w�/�@���������5�lb���ܳ����elV��q%33��;W���D�au�+��UJ��Bn�d�Wd_�wg����I&~)r$˅��&a�M��'��\ f���)`�����JE7^���8��b
le��M��g|!� �3͞�8;��	bx�Fig-��������lw�����I��PB�-1Gl'��F�@+^��U�����\�a(W0�rl��s%\���i��j�e�9���(9΢t���|"�����Kh6����hzҵCK=؟����~(� B�Hf�n��|�,f�Z/���Bڻ���4j�����f�At��p���l��}3#�\�_'�(Wy3�`���ڲ[�W�E��ӎ�����W�鸂Ŵ��FM�f{g54��z����)f"r��j[���oƃ��C�����-!e�ۙ�P[h�9���%�H��6�z��	��@��!�+T����"�Ϳ��(��jD�RF�f�1{Ơ^b׸g��%ȁe�+�ć���Y	�s�;�������I.��jq]>��{�B��	��_-��P��1s���E�HNx*�"��	Z���R�Rj�Gh9�^++r&0������:$c}AO4�{v��\b��==�O��o���Ԡ�)ᨓt��#�\♍��Ѝ�$Ӕ07�m��J�	�b����"2�H�#@1�0k񴣼��{���z.;�K�8-��:�Ԁܱ8h�&*N�'|��4���?�����h��9�͔���sk:�V;�����z����.V	베ۏ-�D�dūk�5ވ,P�Q`-俴�P��ո+P�}�jͶ�����e8�I�<{@�xJxנ�|��g-�H7����x���<SYB�%���A����c�,���Ǭ�8�V�2���+l !����U��U;�+��eB��i+d���=���]�PMe�ML��퟾�j�O��x[�z�;g�������y�kƌZ�*���}�kP�G���@uO�^қ
�	�QI�~:6����-qwqW����;��`��Ќ�g��忛����;��F���Z�q�6��o�J��b�I=N�.�p��v���XS��=��??^��ޠb���S<��,W�Y��Bx�E����b��0|������E�L�j+��Ή[t%�i����~A����Q}��?��1�6��� D���\��K�I�®E��B�{�(xaJU��D��-K��*'��~�����J~{���Ҷ����#1�p�M�������=u#�$�	��
����|��֝�ۇ���fy�=����}��.p�i-:J��P�� �H�FO�A ����\U6���06y���_�F����.��̎/�X�re�?%.��xm�����[�}���ڣI�f�&ޱi�zLz��o�X.P_Z�ĥ�ۓ`�=����������x�RkK��" :"�'z+��m��R_0�H�=\����g���FTB���8��w���:n�pxe�y��M���{�[O鄽�
��oU��0�PƩ�2�?�SJ���+�ɮ=����%]%�ʌd����7���?��0��-@�Y��1Q`��Щ����� �����SgP�-7R�]�+��d��퐊��:��Ӵ�����1���-^�XP��/�vǒ���涞_�ťW��5Ӝ�e�(�� Vɦ,�Clw�Ԑ��Sfp��zVM�Os� $�d��6�dd�P�� �B: !���$=��ϯ��f/#��l���HO�(��<�,�q�sz����ۙ->��u]�Z�v�^�����S�����}�~YI��s'(.�;33��h9vz��d��iuQS���/0�����$4r\�M^
�ݚ��xE4��ݬ��f��5� [����#~-�b�MP������r�_���d�jeLJ�=����= ����a;����m5	ܐ	��e]Α1Z��W?ֹ�F�k�^��_���!����Ԥ�#��c�K�
�ZR���̚���1o�o���KP���U�[�V`��T�i�������e�8�M!� �gxm)�껙���O6����m����~�FڍQ=�Bp��=_��Jk�q|����7�d)^6Y���L�����\;�,��Q]�E�l7�.��h��Wv��:��'��2t�\l��3H��9:��Qk���Ù����I8�?�@�g������eHi0��ڝ���?�$J+
���{�m���N�Q���	FN�2'�����dq�Gwd�rZ�
�w�@��?Ű�Ⱥ��>)��?3ڈy��/o!-"�Z�bַ���vD��P��ܨ}�3]HB�6�7�L������7�N�f�u$R����'�u���e윺��U��Ty����x~-y?�q���F�D��x!x�.yUIgw��S���rL�������8��ߛ�U��/Z#�p".	-~�qJ�S���ݧ�R�Uղ>'/6������c��m3��q�R�����]�F*�Ķ�M���Q�qG�l�a&j�[�\�����;x��7��9��3)��'�����M��|�G?%(�WM�W��ۄ9u��dot�n��ϙ?<���i�8O �_ ���k��ܵ״/����z6f%o��SG,��J�BU�����,E�zP���dvv��!8����
�;qB#�BÉ�2����p�)8�&��<��D��L�����0h��w_0�=r�����.��A&9�O���k�l���<{{��G��z�({����A#���U��"�[#��m]��^ ���X�XB�$w�/W2GydIi+�b/��"�Y +����vO]?ɀ�B�G$<B�Љ
ad�]�Խ���Sp礵Y���Ms���7�\_'�rs�%�	;�YE�,ԑl�;�(�J�����k�+����{�p�\���3�pa%ơee)�75��p�����"߳���69��}ʵCM�q���λ��i��%+O6��@SfnH�1�Vv*�%f��?|�\A2�QD�7gq Lc�9_5�8��ў'D'^QEGm�hUU{�'����%��WX��aR���6�d�1�T+ [7یj�N�P(���q��'��aj>=�@W4�4`嫝���DntBn)�{)�G�T}�		p���q��m���M~� �w9��~��B�X_9�?|�#�fφn��/��o�.f{���t�ǥ�Eă;�@�'��<9�6�c��3��?-U�!G��x+��*��h/R#I��\;c�1�]sU{�ӗ��*�/.aQ��Y�qf�8��]I7�Y�p��Dť�T	hI7����h��_F�7�|�Z��(24��+��e�A��,�,It��P����n��l(��W^��l�aǋV"d���v?.���1��J б����3��maR��?	�������*��Tb5T�C����rE����5t-�"�:��!�W& %��7�o��>hj@rK�Ѣ������ 
D�1Cz	��������=�k��7�'BH{�O�`9ၤ��0�gW6�j�j�&�M�P��VU+���ջ+0l#��^3OD8����?ԎdW׊����p�B.��� 8�����C�u:�:v��{�xb�Z\��L{�u��Ss&ڰ�1��)�ㆄ$����{�%=�=�XL)�T�NcK@K�VY�#{�3� �H7����s���r!�Fܳ�_�����TA��Uh�`0�q����@ �d�]���t;�hVE>7‪V:,�J����X#]=3B��ݣ�� xZ��"D�r������G�~o	�(�A]��u�~g�/p���r$OP��z�e!���-p#5ò<�e�Ru�����Nզd���,�1`7�D)^�Jz��e��;mv?��n�$�W���H��t�jFzQ ӯ�yYHn��,{�r�,��0�^Wk����a�g={a�?���J���Hh�ƏƜ��D�T=�j��i@�_� z�R�2d�yгI��N�pg}s\N�����������6����
�f�@�R7����9�Fpz.��^�� ���Z@�s�l��=��]�~1P0O��,H�hC8F��=!R��|��h�`�0�:�z��oZ<u�o������	�xxܩЅ�8�=T1�6�/���i�<��4�1�� �<�cw�;��������	��朇 3i��0�l��%ܼ�>KgJ�;l�g�HQ�eT�� �(�U���Aám!د'�/#��,�������Dp�9���CAf;3K��RN�N��;��Pٽ>�HU�7�F"ڗ�j���q�<pj7oi)�r�{���t���؁d�N���`ɞ��c�y��"�8*=ŀY쾴��"̍r���C��Y�� ���૊5�-R�0Ϧh���uKzt�c�+d���"��	U�j��],%t�30h{�奚�ۉ�H�N����� �i����~!
�Q%}�r�,�k�V}"��L6vW!	�����vH�ދTB?�n]��~�'��n��WY��ev��I��rYD��)�'������4��+Ѣv��Q_�>�UH4�g-��趧����r;#`_�0�����(�-�ƾ��k�q��Q#u�λ/X���C9���J���OO�h"�1t��ȕ���he'� �)b�'j7h~5WTaR,s9�K^Ѡ���O՛:&�Qr��'dPβ7�g�th�IL����߉fwu^,L���0k��A6.�$`�X�qJ�	ѱ��3h�}��֌�:gLYͨ�@r��h�7��1��9�s� �<���#�z3��^E���Ϲ�?�#)*ղ�P[��A5��ز(��{ć���׾�D|GY��l���H|哹�_��b|6}=�)6pɠ�� �VV�9a��Ń��+߄�^�S:E&���Mۤy�eFZ1�MISsѬ��Qfէ�����͓4^��u��6*fQ�s��e{l�Hn�'�����(A�Zv�թ �fPM_�EJ�"b[��\�MS�7�)���k�r��Z[_�r��~w(�	{۩+
���癱iZj�: n��16 ��l֠�9�0au�|(:��m�Wk�sU�����7����۠��E�J:Z��8I:�&��=9c��@��/pHa��6�&��~�>G����ᒥ�@tR���*�-Ń�)ӽή ���_��W��k�D��cam���Dc�<�k�����	 �o�����0U@D�\��3\^O�Iwv�1�Q����A��sVv��XTM���P+�`��LD�m���I�%��bv��TM�����������hi��HLdM��FieU�+��h����hR�s�[A/*S��O�TP����=�H�躭<�������ȶ��?s���9$diǯ6l��k߈Ml/�
)묶�3x��QLP�F�"}�8?s�U��20S/�p��\�^���q8����mƮ��	�$<�}F��N@��pE��C��TN]��2w���a��h�TeJ�M]�_-*�Fk�4KKSܼ�����W�9��N�eQ����cķ"�%��L�����%���%��;�猦�<.�!���	bij�c��`��}��%I���z;X���PȄ�l|��̻G=Q 3q�o��P@h�|�7�pb������+�߹<�i�������=;�ފ���S׵�l�v��B��+@��`��x��{��o������n�J�%��fyp(D7CC���e!�o�'��w�Z�A�'�
��0��PK��?�&\=�r�aZU�o�@�/�n�E�E�� ����|J@�W�]x�JC��{ў��7�҄���P�2��j�m�bw*���ya�o�E��%	��G۲񘥥W�f�KYU��0}7F��jQ^�%�[��Tg.�����O2��9�-���9vS�Ts1^�Kv��6��Y�����{,�Ym)j������$.�*�.�b4��Q)c{o��'�pgީ4��۱��F��PT{n-��'��h�=*o����N�q���GK�m����ɲ�,I8����'R�J��3{�Op�� f�@��(�wgy[�Q�? �H��0�)�-�m`��p@�g��Tu�U��=����G��5�[��`ц���A '��`<�0��e�J\,�^��ՑY#5砧el��!�-�����H⣣�(��!r�^o��x��{"�Xj�-�����=�M	>E���%��\=u���R�{0�$L,��bGnT��A6փt���ⱆ.�<�|],w��Q��o8��P�\pa�Q&c�ph�`�c"��9N3�eS��@U}�B���r��]���I*T�~����P�wwT��ɷaz��x}�,f��E���[#B�N�:Q�/x�꾻��R��^�W�uu.��]�k�.f=�][�z�"zw`�i�d?0����=��1��^5E�G[���\)P�^�A�]���Ktx�(�v�GU9�^�q�ݦܔ���=��k�κ�O�x{�<����Q������j�J:��(fH�U�;T)=R�m�u>L��ֳ����C:*��CM83eN�/�\��Ծzt����X���w�xTS�D3�����S��-[R��{+��Ph�r,�t��&
Pc�,s�պ�*��5?�0_���~���������g.ծ�������2l�f�0E}|��%�a�?Z(�V�I����8�b��\�a}Tl�|*׳��}\��ɫ�!�j�
����\��I�U�2Z�@���G�����ۊQW��da�n�s�1���{r���6�;:��{��͛)_$eN�i���ɪ�.$-�HgW��WB@�O�Yzvm~󷃼Z%���զzr�J�F1 p�����ĕ����o�~����VfsI��?T2��%���2�ߛͩ��d�7Z3��rc>�`�K?�o7�ęl�Ϥ��)h�ìiJ����%�ߥJ���H0�x�6������j�
�l�tW��ю��S����q���_���g]��\?�t�>���_�ݾ��=@@L.e����(8.4�� �?x�L���VM��j�����T��:QsХ���bDS5[��� �R[hX�YK��$�t"��9�q)��	/Xl�fŚhaoNe���	�dD�����<OwT��������3��~h�L,ް�
FA}&�H�S3Y��;� ��!�Y��pZ�L��VIR� ʘﺞ!������s�����"�|P�2��>�($&��y�ĕ�Fj�/s��U2ٴ�ND��I�O~���|6��D�X�1��+% �9���T�������؞��01����ك��[+C֓���?4$=��&z�\x:/�c"ݰC�%�����%p?Hd���Z�
��W8��C��{w!h��4/���:���<jWK�/��8��M����I�H��QF)�U�3G��]�7s��Y4,ٷ��d�5-T�ݪ9H�K',_P+���Ս϶�������E�LϏR`�"q�V��F�� ���ݸ�>ݖr�r
�J�iW����7��& k(�x%�C1�����A;y?ݴF)���� I�I�)w3Q
ȩ-�l�R�G�`���PnU�&��f�m�f�D��H/k�k�DT�����U�"2�,BL� ����Oyh��Y %|�AΊf�[p�y�庨�2�����,�!~�%	�#�-��U�ƃZ��U\K˼m��J��"�8S+2*H��N�됫 J��ݿ�b�Αԇ9�3��X}�3���D�e�m��6�[�-����6R1�h~E5�
���B��o�V���h򖺏!L�Aa]��s>��[�%c�Z��f�����V��J.�b+L��qzT�J�ў{�ƍ�*'/��G�"$3�zm�v�d�m��i��&'D��)���e�l��E/��Y�t����	�աȰ-1u�d
�t��7�F�K;���`�����e#�@���U�D��h��RO�
�Q��e����y�]|+�+����!+�n{����Ҫ��mB��.��A	Ns�"A�_�L�e�Df�������3�<f;��F?�� �L$U܀�81
u����16����/�&Q�5�f ո����mcY~L��t \�Gx�t}e�~�U�N0���m�(Y����Y֛^��G�E?������?��|�{�9�Ѹ�p�`|	��9�RGd*?K���S?ɗa��8I큈�g5��2#�T��� !M�����tT���'P.���9����8�0g�u[
���`��2�WLwYZ�am[1W�W��tY'�MT�X6&UeN���E[A� ���d�q�U�k��r��˒Br�o�%�"H8��4�$�`e��8nL2��>�	qϓ`��%:vI=e8�(A�Ɲ���9����L�9���k�VE�nZ��F�q|M9�X[V�ER"7T���:�z�/I"(�pLM)��,��1���QÜ A��(/}?�ڼݨ�e�ϧax��lV"�9�.̕Vm�́$��.�����Q�g�xtR��>�u���+g����q�CK�N�uڔshg���ާ�(�yKB�E��+A��%=�F��tȄ�Pj���
��b��J��޾����.I��;[Eh@U�y�쎊�ET�[V`y�F��ALn}����e��_*]d�2��1Yֶ���q����[ �̂:����:�_MY'/vC	�����௙V~�~�Bo�Щ�G��+߶��MK�#�?���K�'����[t~��Ŭ��k�>C���p���ǭ
9�W�웅��V��`�"�O���Ϲ�<w��拷��)�st�ݗ��WE�C�� 6�� �r
s��3� ���A��P�6��Wjh��E"w��rLr�5�YeX�P���g/N��J�]��J�Y�u?C7��I=p_8��9�ʚi���xq�Kg���j��TS���H��Y���H�K� /g��Pr�̺���y,�F|�L%>$"�pZ�Oz���g$�ӞO<N��КF1�G�bj2)!^�.3��X�[�l�Bw=�X_T��(_�#��Ţdn��ҫkIUN��eXPdW��.�}{����J�+�7�޳�U&����L��"�3{
�G��{���F����1�)���]��%����s^C�n�$Z��i��IY�=�0���	,4�(X4�wR.�U��k+�J��"�����m/��y0>�owL�����jrmhJWо��;&��C#'��5�����`�����>#N������z8x2&�F�d��k�C�����Z{&�S�h昭bQ�
�PU�?*�]<{L5�	Cڛ��8��7�>v������|�^a�aU��A5vME��=и�BPO=�4&�W��Ft�-w�ÔI�U��"L������杂v�B���oQ,,��	3��S��ǚu�--�I��AS2�k��iʅƆ@�:�"3�������(Y/RP�d�<b�n�Ôhk��g:HW̪�ڿ���W߉,�#� ���� ���������|q�QDP#��E��i�^N	y�2��v�g<B�LZ+�=T۞��ft���%�;�#�3��sPU��5��i+[��#�T0�*������E�!�?��� 9x�z�1	�d��h@�-���QP���׮Պ]4�?�m�(��u��T�|�����*��u��f���sݯ�C���$Ѳ���*(�NRCE�2׃+�!bJ�뷴\݆��(�>ښ���e+��J� �����GGJ�^��ؖ.<�&��D�����7Ƞ����W������d`F�*(��-i
��ݰ$�#�"@�ܣI��pU6H/bQ��䅵������r(��p
4LZ�������PO�r.���%��� FGloG�D�ˊ^��;�_��wԀ(_��nqu�rD�Y��Ǝ�g���y� �sЫ�nT(&v�0y�-x�Lz�2��S~�14�t7c�M�z��z��1���E�Bb|ˎ�3��Ȣ{u9�$Ydy:�R@��f��x.�ir�/F'�����n�c�ӓr�9����!��I�d�<�<�j��mɟ�֨��ZՂyt��G�/�ܣ8[r�b��kt0��/?#pZ�"�2$	sO[T%̩%Ƶq��~Tq��H��L�;BҌ��U('o$[����G��Y��w,��/��JY��hQ��Ï�¡�2�W�Z��w�2vG�4C��3l���<�?�V�i�,�u3|�*MicsA9J�A+m�o@`6���>�3F�W Q֩�����Km29W[{���\��d��Q�8Fr�$���^U*��i&�h�͕���~�^��yQy�l�!��U6�^e�Th�����T A~粒�4�K��F���u���e��������(�߾R�S{�٦��Y���qۇf�����p���I��mNȧX��ѵf�1o�_C �Q/�F��Ѵv%1	:�B�"�n�E����?��g&V�tܢ
��������$�Qŀ:D�����f��jd���<���3�w�'����Р��P��+0�	��0L��C����.�Y�x_YxAKu�)J�g��Ϟ��o~��_橈f}�c������9��rIɀ�����G�Ow�]���� 6�O~��iW��(��R"��GF�˯�ʪ��K*vN�|@:đ��H���[� ��M 8EJ���Y�V�M&����l���aK���b2�.턾Hk�(G��Y�jn�[�/&����d7��_��S��FX'N��ݧ�"QN�̎ �Zi]��ҭG���%�+��O�-�
H�h����GP���-�/8��L�Wņ���h:^���I����i&�^�S�����-}�j�`�Lɦ��X����n�(ù.��I�Y��"���Ь��9^� �MI�h'2��)�"�Z4 �"�����g��e�Dz�q��3�zE]6��������Ü��l��)�碚��a�]�f�?�H&�9����D�='�T-� �Ȝ�
��Ka|�ǻC�)D�1�$ϡ�%)���~��g��\�tQj�?���+�u*��aF?��-�3ۋ���ix��[#�
��*��k��V����u�ѥ��g`)������R�>=6��n9�F���ya>�(���Ϋ3�����m�)�f/sv��-�7:�*1�ߙڱW���S�C�T}ۼ�7	tf�~c ���X�@x�p6 �Bc}�Msl�G��U����q��22��`a����ՓT̒�w�� �C{��}+��r���[�?�����X���k�ׇ��#4����m�-�T�YE�Ԙ=�]�ȗ"�����y���b:;E$�s�VÁv�V�h�g����1�!*�t�/~��}w��f�⭳�;����;btSo�"<��6�����>3����4���P�N�<��E���d6j%����&��}-�C�`��s}9/�N������$�=���Л҈}����N4.?mt���1^y��@��
޹�F� �"�L4�*
gB�[��*��E��J,��X��9G�d�ޥ�zp�ܢ�p�u^�Cr�T'IFl���bV)_NJs���p3�|Ŧ	�Aª�����K/M��ه`������l�ȈP݌π�p�����vU���6��O�ܶ����P�[�Z�&V,h�����ܳ (=�O�+Ƞڮ�r�z�R��ɧ��B����8Z�ו�p�!��.�n0���Z<�c2Y��]hqo��ޜqck��ڇt��R�?1�| �c���͹��Ӎ�>�(#Ƥ�cIx/�0@e�t�u9�#C�5�?�^���^�MƓ�"�ħS�>��w��/�H[09K���F۞1)��I�D $��j{�~���u�]���w�'���M����q}"�QHߏ;[�ټ�Mw�d��!�A>\B��4�u}$��
����_:�['�C��QJ9'�����L��-c[꾣E�L��?w�n�MG8n�	sc顿���j��G��s�;=FU&�c�2�d/�e�4x!�ga�jڮ�.c�Au:j��1J8Do�K�$�{uK�(�����t�2�d�l[R����_�_�WBx��5�4k��2LG���@�[��E�a��_�Ƈ�r��Αތ��
w 8�]L��T��P����"��F�n'ң�������4~#**-{�B-� +�t����_�-�������1�Ͻm-x~~�H��`?7*1
��m��c�s���}vt,��xgmS1�o�i�{7��Σe%�{�T�Wjn*�g{�e�h3t�.؆>{ȴ�|a���m�������#Ņ�n�~ꬼ�,=X����Ijř#��U̢���%o���1P����gZYĆ*-�;3��LJ��?O�	ݚ��n�p�]�y��H�����݀�r���86�ťYԠ~k~��^js� l�M��'�K��u�l��O�*s�������O��4;���U��csK�֤��Z��X�5w-V�{X�Hx�cL!���8w���PE� :.e��O��u�~���2�Ύ&�q�*�@��߸=�wب�^ݚ)�S�s�Ӡ����ʳB�M:A$��!�rb1���d�}�}�r!�!�@����Hg���I\1�j�G����=�O͑}P�9Gbp��Uaz��x!_�#�xyh���_�s�}��q*"�\}��#}�>|n:�A�\$N��Mid8Fň&���T`b���bH�}�w�{����+&��	@��)*���l�xO=�9N )}���3��@�T��1,���g�>����&�p<E�d�.H1�`*���ύ�xr	�x��=�&"GWȏ7E;����˯�#����)ϣ2���s��|*C����C�i5�����	d aԐ�wyj�86ƃ��/<=�U�;��g�"�'$��q��z���C]8r����������Do�C\@��jLk��N�U����0P2��xi՗����]�n����T��G�{�[9�*������p@o��؇��p�v�8����cZ�A�&�����Sܗnx������TObk�qdYր��!��w��w��*�T�[Ș��u��'>�H*5���W�6TV�#�#��e��}G	�q���/Odg�r8�I�r�Z���*�b�=�M��Tz��?��q`R��o4�
6J��D�����;+:���x@Q��OD��P�;v��J#F��6�R��Դ�x��jM33É�!cLeξ���ѣ�-�ݼ�-�Ok��M���
��JĆӋ�M�RP"�|f�V�f�"f�S���"��-dMq�fGjM@�X��s��8ŝE���1�})��u�L���&�/�������#�]�b�U��|wT(-�2�y#5���q������L�� -�G����#�����{ �n�!=��ԧ���2�Sץ���Y�:+�.���t�^�s�'�B��>iU��~B_a��v�y�W�"���|���9HsC��(7h���N�O7��q�)�f�2�P��(~�I�H/������{�l�/���mK��r<����ɽ� *b�K>��Q���Q�o���t��e�������"��O$�3R�0,�q���)_f��J� �R�j����_�e��C���ݢ	�
��ka�������r�]�uF������C���*1�O�I�H������D�<F -�t��4*�� f�H���pF�g���aԐ����h\����/L�|����#�����/�<���SBkt�L�ok�o 6u�jJ.��x��Ȋ�F�ѣ5��ǫ�.��Q�����Tt�.#�4�*��7Fe�Vp������.�m�i5��{�U�4��d�l�f �ԗ�hO��_��e�������N3�"��$��?D�s��ԯ��u�����4��D�D;�!W�C���7��y_�r�h��>�>Vj�̬q���ᨛ�+:0�P�U@ 'ܞ-3�z�/M;��^Ī��{�TV���1^�K���(~���o_�K8�r"���x�]�R��`�;���ة����K�7�$jO(����zm��TpˁSb	1�==>}L�|��x3�e07��yX@�3����Nd��,'�o`�ɐͱYN vd�{/�{7�0Up��h}q;K������	�</����@��w��\�}��5d'�T��-#�;��El��e2��w �� Sv���J0۾b@g��V��%d�g��&-�6�����۱�	��;���	��q�f�	����X�$���H�y�X�'����0�ݱ�0��,Xc�����G�p��@�ʒ妽(93�X������`���b|آ�����pٗv!sL� �~h�7�f`�/<^�j$'ǆ�
t�
����<��Cx0��<=6��W��íS}�im��[�[1����dy'"�D1�|���!�y�Wi�]^��H�]�f��g_ȾF��L��9Z�C�~x�L�;�/��b���*��"��:�0�'��Pᛊ<N��?�x��\�����m�&���b;(���ٕ���>?P_L������(ICr�|������ףԾ�hNm�������,?��������W���mzh�x�K����BCMܘ�ٔS;��z�E�^�h�ѥRz{�c���T�	�ؚ�}1Ri��(g,׾|�M�(�i��lCP#v9AAD���7<�X$�14��]L��~���i�WH|�zv�R!�h�����������ɿ�~0�Xٰ��	�,�0	��w��aW3=���H%����c�y�H���E|���k�_��Օ,ݗ�������ѝ�9w��G̣	�B����c��~la�J��T�]����[T@r�x���HbEսVxiVr�;��*ޚC��7y�w�I���'n/(c�����u��6xv�gE�ػ�| w���_�/�}���lH�m5�oA���;8VH?��%�����l=ҩ?���:J�' Qm�As�|�C�O����U)h��cŪ���F�1�qZr�o��w)l��f\��� 5et=�q�����hר[��)''H[�.P��$o�����@��@x! �-H��H)���9'�� ��D1���'�i�������:�mCR`X5�R��z�+0�������c��Uw��lz,&��G�hͿ �ne��E����{�A�u7���޽���۔~�F�OЊt�=w��&��c��U�q7?s�L�m��T��r,q�t��S/�:-;p\�S[���Q�\��1�a�s����?fI�_ T��e�;1�Qr�P�
.3��t*�#� ،�F��3I�W�{��t
��WC�/1/w����HW��؆��b�E$C�F���׷�������Ұ�Fx\�㝱�*���Id<�X�bM��J�G�uˢ�U�1�դ�Y�����X�e㷲²yx�s���}D��Q�ūhp�;ܓs,&s� �"�~��_7�|��T6x�L��3.�[�m$�l��-P�r/���+﷫�ٿ���?��78j�J�C�_xyT�P��U/�u;Ƶ1�cob�6wi -X�F]����7�Ҫ'a�;j�p��&%l�ՍsuqxҎ0F�,Ўe�u��Q��t���8��y5#4�;Q�QV��P脽k��R����ʍ΃��%|�@�������u@M�Y�hB�F����h� ~D���d��W����L]y'O''�F�Y����VA{W��� ��-����cB�h�@ə�@Plu���9�"�����O�
�`����Xh��$N�S'��P�X�����Tz��/��8B�����H�bЖ�c>����s�.���f�V�-��NaZ��9�C�9�[l"X$����k=�Fu��e�c�gQ�/���uAd �*����7>P��F��Q�x�a�'�0n���k`�_��4���4�Kj��p�i��eA���
i�ґ�h�oںW��q�tP�Y���(�8���2�U��b[3�cx>��U��k�M�;��0=�~|숪����:/DD�.�5�+��T�Nv������ǲ�|H��.�82(��r�y-�`8�Y�L��s9�YP�6�/�̈����H���	���u�BC=�]��)5���m
�{tܰ2��O��ƨǫ��c���98R�,Di��,��C���ȁtG�31|���o�I��;�,S�Q���E�Z�����	=�����a��κ��
 ��e���!��],����a?H�;g_�ꔖ��2�6��������~��R�Gf]�A�:�WLKom�Hg�����F���I�����VA��G�Z��I��l��>���x�{����W0�cUj�M_����q�$���}$�PYG�V�Çyq�5�<G�9�[�V�X�Tr�7�ٰ�)��4|�S��\*]��24MC�ϐV�9�J	.��:֑�=&0JZ� ����qR�pk�mi�_�%u�7��#�v`B����O%�E{�̦�������ޯ�$��c0�ZIL��'�ck���z�:2a�6c;I�*������,�1�Dq�>r/�]1�+ɞ#�_��ZnN]`=*���K��n�U��d�=�I��R� �9.
O����^/:�Tys�A\��e�{�Ȅ �
����?�0����?�3t�{6��}"BZ��������%NZ��jw�7�{4jU�U�z��M ��6��"G�̀�_���c.>w�5X_����~�(m��5�������%@��F�]P���vA�K�R����ii������^'�O�ʝ���h@������(@E��[1�ݨ��_���D�N,�Үp��9���[ �G��� g
���#�-���ު�}��+��'a�jă��v��EX�l@!IB��l4[��{�+Q��E���hZ�3�nD�z�ܢ�hlVd`S}7�QCF}�tGu�z�;yiVg��\���m�yWn0� r�q���i$�w`��JiO̫�x���Emn@/����F�����D���Y}ц�����9*�6-h���e�����w���/�+��:�n�'��L#��	��W��I@\Sr8��*�P}��^��7Tk����Js��\tN(�̟v'��W�Ȅ��
�r�To1_�Hxf�ԣ^+P+ACT�4Ds3[\te��I��.���XlDe��M}���0u�2Xm!"�KC�Qc�W:�ʾ|���󻮌�{D6�+XxAډ�$� U�ɐ�b�	�_��I4�y Dy��tP��F��������@&��f�WURC���f��4�����c)�#ph�{9��n������j~�e��|>�9/�
�IcE�/��C��-X�O��{�h�7d�B9�t]YsB?�)���ȕ��˿e��6���@���r��f0�6�U�?H��G�E0� �H:]>{�@~u�p�a_���_H����0��ZgX/�Z�Ű/e�]�������A�W�S�bޔ���]���N	o]��[��F+ <�ݧv*s2��4��L哉�o���N@8
1YRx��a��#Rj���	≺Mq���l�#��oH��C<ud���zU��DäV3���N$�E�����,�Mo�E�B���V���/�o�$>�I'ne��U%z���������ż��yt[�������f��i꒩���,]�we�!|TՏgt�������K�FdY��wH%M�����fG�#B:z�⣢�Ҳ���O�o�D���6v�V�I�aB8,B`̬e�P�<ϔ_J��D����ߵMhw��f!Z�*�DفG�Xw�GG � �#1c*��l��Ϝ��A�u@\t7u靋:����Z���<���_+q��&$��7�B�f��k�&���]+��Ѱ�Q_AN}�q�&�l.�:���Y[�R���#��U'���|a��|�D��A��������#[��0���5�K4�"9�	��up��ҙP�JJΣ��J�H���?_B�Wk�؊>�Bh�/)Q��������>N�=�m�3��S�*�J(�Ҽ�E��Q���	��"�r��d7 -��e�v��ޤ"�M���tI�i~0�<�ٟ���}���nX	��ɂÊ�+����LH���R�q��� �e��h	�C_H$y���ϳ儩�Q�D��վ\�1��ua��|�WC�@��^�{W@��zf��ۑXZ���J��&c��� ���Xޚ �dP���@����@o,�1��uZm�O�ŧ�lAB(Y����R��۝\we���H�SX٧у_�&2�/�<�q~|�o&N���^��ҟkU3�ќ
�;[WY*���|Y�:w�g�Vy@>�M���l\#II�=eqpX��B�N��=�O8����I����d���%�:���0&)Q��|�W�5 ��%��1Լ;���9�����+�(����G䍾�I��5��P�O-�Z���(�Q���Pr��pZ�����TV���g)�/��������\��£x�A���h���pWL?��m���=V�r7�>e�yT�ؙX�C�3:C~��ڳj���ZQ=�u�5X�|If�t0����Ŭ��|�cJu�įEz����a��������h9��Л��tWۖ�DթY0����I���֖���7L��,-@����O�)� �qt�1����c����m��݃a{�9����[�r)�,�����s�!%�D�P��ͨU�B0�͏)
1u�J�T	ٸ�߻���r��Z��I�PP��zp��h��/�N}�@Q�c�M{+��w��~v)Q���Ā�eӧ�u*�y.���@�6�K��ᚕ�ڛ�*�D'�v���ԅ#ǖ��8���'U��ˈ�������ܓ��V׻��֜���N[l7�WospYȶ2��l��΀�R�Y�W�AL�* �>L�N�8X��YtXf.�i
�� � ���*:�����{�R}���č�gU1S�;������U�ViTnf�q]���l�d����Z���x�Λt�r����eb�����v�����Zgk��g�.�y_31@��H���£��/��J*UD���[�}D������ֆ�"�%5��s+n?�m�0�Ƽkn�c3���E��&<WnA;��	����
� byb֣��vIP�0]4���5���&�N<�J߰��Qv��/�;��;i�̊�H�ᏂS��5���{��M߶h�E�Y�.��|(fR��kb�c���'�X)��F��N�5^U�oLH*�h���Zi�ܹ" M�`�~x��}���2�r̎Be����BeOpy�}�d�p��S��sU"9V^K+�^�ܘ������s,*C�or�LX�vlJ�n�MV�h1C��� �u�m�n����I��z>�T��Q�0�\�^~j���]�� ��싩Gk�F9'������C����;!RT�0V=G��Q����xc3�a�5,
�����&ċO"8xyF9JJF)��J��.�Ө;V1��-}k'l	�H�KY¯�Ta=�5;O+���?�
q ���b��o�����Pa�C/�K��y�U��k1W#�	�j��v�� �b�ہNuoE����H����v��ؙ(�]*G���J�Em�'�������/��e{uFi8m����ˮ�i��˴k��v�G�D9}�����EOLc��z��ƙ
����áOߜg֖V8�l͛����q�,i�a�Ďnp3���}S�y.�"O�\U�I	���{���e���V�ca���#;�F�`���Q�O�)��H�MVJ�i;8�V��0��K����O����G Ze{)Ձ�W;����T�v+<�-$l.6�7�ARA�&*X�0�S'��c��)��A�ݱ�l�,�����D�O�>K�e��8^�-^XxT�2bw�}CaQ��xZ3�Tݽ.ۊ�>Ƴ�ZDY��:�?�D-���J)k<��Z��'��#�ߟL�5��q�-7���l�9��,ܠV$�+{Fî9�9�/�@��ٍ��{X"澡�,��@�@���'-�7�xe��������6��h��i�\qn��f'�_{��	��xP��[��Ӄ2��P�Z?֌�
�F-w�>��,V�/�i8V*J_[g�v�";?�R5K4i�TI��/	ĝ��դ �BP���w�<�*�8љ�{>_�^��u�OC,�
���<"7az�**xf ��y0`�Ђ��j���X����6�0��z ���h�����*e�����u�@��N��ߢa!(,惎Z^$O.�FW\�F����Մ�$g�}�/�k�VbW����V�MN������a��Y��QGE�5�݀|Qk�� ��)���V�W��>�R���us�>��=M`\P\�8B���v|��I�V�"��:�c2��3>S����q|�}��XSBb��A�M���4~�/O*�x�X!zr��j��oh*��C]�����~�=9=��X��ɮ��|�h�������W��@W�ipve���ӑ���ݾ�VF��2Xdf���ȯ�RS��Q��Ƀ[
���c.:�}R�. �?�	v���:$�4EJ|盜�%]�(һҭLyG[p��2�`����π�e+� ���@/����g����������.q����c�Z"�XτR��O���b�I����2�ǀY�BnL�8�e$).�j�A����d�3:+���⬚��Q�w��jo�Ti(�!����d�Qc,��ZN(��Q�G�K?��1��� �cl7?�-�ni�����2��	8�s7i�gۦ�U����
o��/�CIb��OD�u��>��1�P�wkw�ȧ�wZ���ۓ�#��S�"����s�y��/�x�0�Owð;��ڧ\���Fz��s� /S,e���N��x@RюECc�r`�k&Ahh��#	Yw=Q�zD�MGH=�%��K��Tj�s�v?+��҄�����]�9��-R3�}�*�o�T���q�󤋦����Y�Dp�h՜6V��{^=	��5J�l�M�/6�`�\��P�3�Ղ -���Q���C�1�}�ht� �h�)�b�95� �!3�Z}��EZ�:c*p�ol�&��N	��UT��������/�~UoJ�?l-9<��=��cx�u�)a��H��m�����ܰm-��Ӷ�o��a>
T�UkVX��^�$3���ɱ��^��E�����f��s?m/�Y����Edtj����q�0���{q�O=��W�J��7���	CO�h��B�qx#�t�������cs���l!PVD�ёU�u	OjC��H~�J�tJkd���	�߇��L�_Tm"�@jBR��#˖h�+c�[���8)���FMrc<�N�sy��܈߉:��9��x��bղ蘍��J%���L�k���'R3v��q�����������n��RM�t
p��a��d�����L���%$r�����M����V$����� �;$�+������
�� s!m��	�1���[����J\QtxN�5֨�k?��z
vm��f
��w�=�i��#g�0��ok��UV��2�ٰ���M���;(�T�Qu���E�K����X�.��~��.uQ(0��*	D�� +�;z�ݯ,�헻�m�`ѱA�`�0�6gH���m����x�����QJ"ƽ�a0>���зa� Hk�Z��4�}�s�{�r�f�D]C���~���=Δ�j�!�jMm�����,QQhցYCbH���A�W`��nC�ɉ��يW�=L��J���J���1eV�0s!�£J�?�f����8:����~��@g_ ��p�m�8��|&��X��A>�tA�6^��I�{4�]�(�R'�l�s�ZB�iH��	`�#��O�a��#݂U���s�������~���oX�qy��Po�P�g#����\�`$J�P�j���u��e�Х�-�YF�9����
�͐��J��2�;!���Y;��ξ�MZ�n�W�jCǖ�^6c�2��������>��Ŷ.��[_�l���֊�{/��d�x��&7@�F�V ��p�h_�6�*��#,�ydF���-o�H����jJ�oZ����!)��7��)��_�!a�-���6;ʜ�ſ��X��4�����YA��*խ�k��c�vdc��O^˨�U9ϳ��v���:�����do��ƫt�'�x��������J6]�j�,K�pe�#>N�>�i�P΢� ]ͣd��cF	�s'��n�wv@q#B�B@Us��jY���(������^<Ӿ�dB髙�yOaFx�ds�*d=����cF1�P.��~��_�F��2ϥ@{��� #��Ұ�_ce�~C÷���^8���K��^�
U��҇����3'B�ˈ2T�!d������`�KO�)���Sˑ�u�H�b `�x��_ďS��n�������� Z4�,�$<��:#:'\���J�<��#���q��{�<��JL�ݗ�$��ӧc_�y�Qn��b;�����Ү�L�􇽇��Ά���=�/_r�cM,B�dRq)pg{�Ѽ��_'k!'r��uξg�n!#M����I�tp������x!����8.R{�&);����0�nFPȂ�5����o�6���]�Yk�)^��18�=��/|R
��(���N�o�~4��x9�u���~�_������]I��¹�]�I�� !��y���PD�x�AB�ML��m�bh��N����A*���^�;��l�*Ua�����[h%�P��.���B�d�)j�a�ơ`
��ڟ݇���zf/����� ��\1&�-���vl�ͽl'��Y�)�� �54+sq�T"��\W3�Zmۦm��;i%n+���np8y�U�n�»z���l�Nx�§�O�Kϕ�X���-6-s�0��Np2Ui������5�X����̲砘�"�?�=Q�T�^�^>0�T�� P�L%������HaQ����8H����3y&��ڭ�������y����ZKקc�˶�%�a����)%�
�*�`�%%���Χ	Sț�f���m��$���D��wY%�F�%S�qv�:���;��o�6�T�؁�~����,���0 }��.Jx<a�ͤ���w�V�V2���@����9__38j��O����-�%ݷ��:� ��q��W�|1��#���
�J2�Kr�g����:r��m�:N�C
�44-�v�-�dT�9�M-{y��ݭ�Wiu�R�].>Q�v{���3^On5D< �3�t��o�S��w�y���V[�`����
e�ZU�0ފT���O��>����ʖ�91K@An�<|.�8㜃�"D
�=�d��cK�~ �M��0�.���|�F����$�c�^�:1�^ک���,UY��(K�7���#Ȯ�V���5��+�2��"OY�
��	�~�BW�DS��aZ��<�s���$Wj�ʠ�+�7�҆_��`=H�'j���6�i!.�z���Ǽ�C%5M�A��6A�or�a)�R���ĢF���^EyN2U7��H��#��A���HiD�9&_���Ia.�֘�l�D���i����8F���KT^L��ڰ*��=��+��s v,d8.��o��Ɉs7�3�3]��*#�|�̫65��ZyXx������}�J~9
N[Rm�J����eR���` ��޷�udV���P��%`"���`����04XP3���ц�λ)#�%t���L��U�Z���9ҫ �@�JŌ��&��ڃٕ����
�F�ɐ��O���JE��	z�Z�`
�}�ςN�3�#U��ƛ�,�<7 7�ҕfk"�
ٲ~¨�b���X꠭<��5����t��.Z9��B�233��3����n�mU�b�H{������D��Q�e���z���\u��Ӣ߫�X��B�iQ�+H��,��8(fwM!9��2�J��?a���~��r�|i��OW�+~u��T��)��O�c�9���G�p��E� ���2�
�I�U��mS� @�7>6kV��H�&dd�=q��G���rĪ�;=���]2A �F]���X�;���p�=�-F^>*A��'>�����(\���F3�c�3H�� ��!�~ϕ@�3P�
��^��Wu��hϋGܗ�	%�^%>zq�D�l��ve�S��N�$_QDtx*iJ>�M8�TE4�/^r�>8�̫��<rh�0sܢeu�ubF��
(������5USϬ�p��BR�Ƕ1�뢍����4��5�4εd�tLԋ:���gqv�Q�QN�Iu�D� "x7Y=��NZ�kr�N���W�u�1��Gz��3�Ji�3�ΰ��Xw��ɡ��/etI{�ų��
��������g5FeG	:��+
�3JW��G?Pp$��҃u�ݿ��s.bLs������g�=@�g>N���L�acX,��=~�ɇ��e|\�e�
<�򼉳F�tu�d��Mk����*	���B>�Y�����˲��T��2����k�-�4���`����X\�ro�5ʶy:������񃲉��� � `�o<G�t����+�Y�����f<�r7w鯎�Ӭ�F��S��j��qEi�N��R��H
�B�?�]���	dl��&m�4L�������;O���tŨWe2��(xC��b U���@A�vǢD�;� ����\���7���RS2u�8�Q��1���!�s}�lZ�S��j�]�P����"��TI<�4�=�="<�M QV �#�5se#$��[(Ө�S�)��xv@�\��w7����k�/����Ύ?�mQ���z���n+����u�|t��IkX�o�-]uC�	v�
O\k�2l�����w�b %]��9�eA��3��i}-��L�ƫy^�?N�I����_="��^�	�S.��ُK��</�1�3r10�K�c�Ll�����'�
ww��>Y�o+�U�K�4�Y)�)v#�����X���S�0X�tLj����.�H���޹>E�,�R�	5�n�&7�kIk�l�O�2Ǽ�VwapJ�Һ���Kn�/|��َ��
��7`ގFR��O#�΂��J�Cp��Z#~�O��y��1eןf٬t��?�J�v}�u%��J
�6�Ϝ�Bo(X����h��qL���o�V��I�mQ]b1Dv̴���	V��j�
��0���Σ6ڌ��yj��(=���b_����%"3h�D�$=d���;_*���ʾ�uA8��V.�kQ�9o~+Oٍ;^d~��	uoo��=8Mj���Cނ|LJd����E�
C�����Ei=��
�����3�+J�-���������#)��
䛲iKԱ�!Q���Ð�Xa��S�_:��S�7p>�t�D�A�O2�~��M�0��[��3=��N��"��N��"�� �*Lɵ6D%R+ɿ��T]�Kf���%��Ws�2Z?�m���ӨS�U�{�N���-��������fN��Hӌv�	�y�K�jA>B��� %67t�l=j����zz��i�O��bm��C43�����W~I�i��	b�%3�
,p�����EK�Ic�ʃ�����k��z�Fztޓ<�ޠ!&F�*��ߐ��@���9�бwߺ`W����9�u��ǇA>�*Nn&I*�o�\,v���v}lR�ťKY޼����lm�ب�� �5;q��a"8�Ȟ�_Ji@<�f�
,:�����)!)��O��'��u��k�yB*����Y��@kW�\i%U�>AJڿ㈠�Υ�C�6_�\)xG�տ���%8���@��p��D%�6�2�0a�=E5�A#nMk��r�+NA�n���0�&�PX��2��NOh��-�*=�U��G�_ou��5T�s���VR�P�'�,�$�*sFR<�=�l��$/|�d�������4�Y.H����Ң��oE��y�i0֔�M�:]���Б�lp6,��s��J�3�T��>@]��ԕ���=f��-�˅�LAu»�T7ӫ�I���M���� [gb��c���?���W�
��`�s{T��ou8�y7&�K:8Y����-W��B�q�i���o"��5�M�H7s{�B��ފ�0'u+��5h�t�x��O������bl(��WMЖT�R������I���6&�l�O-h���;�N6��5�'=�+��/v�������6��-{��uc��饤at�<,�sc8�Sf(�o梕v�sz^����W���_d����>�kG��T.�JP�/Z{2���A�s�4�- u�F�� );��M2�L���@���pw��H^����gEV���{�����xܶ!��R�&8���8����h"-�KV�_�LD[��0���4�m��uB�k����`Z!���sS��\�H��l�#Z�xT�ؗ`��~+��I� M��0��o�z;pW��I��Hz��
��K�ֺ�y��楢||8YE7�Nh�yY sc����@M-U�bO��~^H�����Y�h�yb\f�RԾɴ�?7����QX��0�<X�n��O?6��_�����Vb���:��u��	�,��H뱏�#"ejH8˼��O��N�4�[�� 7I�FCo�UA�n�[X��u��ʙeY���*֔�ࢬ����ƴ�'�Ec�a�LƜ�UƑ���˝��} A�.d��XZ܎� !r�z�*0-SZ��H��(��Ss;��?�fsu��S����qݦ�.l ����G��GN��!I�*����m�hK�y�X7)4a=��}Lۿz����<�U�ijq=�B1���S��3�J��v�f��M���L�|52� ��-;�~���q\�u©I�m�%w�!���3$9��7�v�7N�����^T�?���ExV�e�u]:�јb�mU|LK4��݌1��i]x��G?}��������<<TDY0�/�vD�Jg#H�M��^�)@�^�l˃�QФZ���U��wV �1X�j2� *7��mp��a�SW�U�s�ڙ�	�l�5 ��z�^p�Pt�؂񲿩Ӑ�:�����2MxM�,9��p����ˢ.s�$�S*�,x�ml��x܇�>'�����gԸ"HA��^�oqs�t�@�ɳD~��J�wAe���N^�4�$�y?\`�E]��K\�I���Vt؟b��_ԎA�{�L+��k
�9���@�r*��ojãeRӁ*m&��j����O�������ؕ:jYw0�>���ޢVp���y.�i_�e�2H������Wˈk��_
J[��O�{�T���J���eEd�V�lQE�6��t�!z)=wX�GA|��!�w(��q��D��2�7b�8�!�>k���ը�F���*���D�f-�qR����_��8'����n�Z��>���<����G()��^�5&S�P�e
�-��^ߤ�n���ٞ�-��jC�$<����Ғ����قޜ��������ҷ�2�P�t�P�Y�;��h��A�$Ms�w��ȕl�d�'�߈P�%w���&���Sjw������PyQ�rT>Һ2���a�З^L L�"��(�u�9� �+����藽f�\�%�?��X[n'�q|� ��4��P�p2���vx%�<��O�<�V��_2(=�5���x��y��`���O�g2:�>W�p���_xF���JA�O�ru,��U_���#Z�E��������L�7��eS��4�ꊡ2���T�gU^�����R�U#����e4`�s U�G�G����H�7~��:��0���½S#Yڵ�k�EŐ�T#� �T�[m2���f�"p��Ҵ�{ )5V��[�5�<�����x-z\E9bq\A�:�݄�a;zkN+�"Np�q�mk1O�G$a�A��ݑ����ae]oQc��2	*��vSX�kVMgF��_C��I�% �*F�Uk�z��5z�ۿo�L�@��씷_��}a ���c����L�;N�yk˷�2;L�<��?��*oqK�6��Ba]���V4|��n��+����o��> �?����ehwɋ��[
=���/6	JwW���[���O%E�x�q�#[ƒ?~G��$��F3��)}��ީV�\�+ưzK����1���3�Hų��tM��G�껍p�4��my��O6�D0;��%Qu+fh�@�]+�|�C��?T_WU��5���rb�]���bGOHj5��<>c����Wi�6���R+�P3��젽�r��E�8Ge�����"&�}��U'\���9�-u�hX�'�`=�3�L��M�,�����Ij�NN�g51T���8M��T_V�c�y�Z^ʵ%��:t�;S�&�g�ױ�!vX�4������>�m� ����\�K%:Ǣ�ܞ͏��Q"��+/@��&����Cz�FTA���-#�E/Ja1##���i�H ɏ���?� �V2���a�X��bS�Z����VQ��w��D�(G�#TN�@�a>?��^7=��_�Ja2T-L�Ƹ���z<p����o�9οT
�\V���{#�v��[w���I��*C�,�)N��Uܰ���U������H�ǻ-�t�m�0h����`��G�:H��Hn���y�6�At��YL�~� ������i�t���xj��?�����O|�k+U���$�"��o�F�j-W�m.��`��Ŵ�C�,
=�x�CR���h�����"1:�,��o�ͺ���z-dJ�y�.��D�9�8oA=��F�y�Lp�S�^N��z.Xi�8����񆠽^H��߯y���'���$R^Ka���P�����a�,6.E��QҰ���:z��]�]�9�	�D5̕`��a]�X����`���=����T^Ϊu��FR�7w��en�/��=2`�/A��t�ߦ��0�wr�`��u�y����A
ç8w`�,�]�$Od����ޚ�0�Uױ��
�[ϫ�m�E�m`�C�؀��L%C��])��Q����+=�{���p���M��嗩��	N�\����$���+���{��1��1(�	�s� �Ļ�D�XL��C�@�.XTf��5I<�/�[4W㟃�Rm9}2�{�5)k���a�Y1��������c';�5��Bc���I���~�<z�ߖ(�n�W襄�.�m�~ �c�˰}�ۍ])O�h�R<�qG$\��F ���9�F̲�iS�yy?�q������D��|/[II�{�n�h��7��Ȩ%�2���[��Ǧm(H!���Y`6�k}>�;jW�'����$�� ��NV$3����ܑ�W%�T���@�5��~����t�\hO�ͳ�T�J�/��<�n?�J
c��
��#��(��r�8�M`k��"H�VJ����f��&��9dl̵�E�_pI 
��	z����2��;y:���py�?�<�J��fw�/�՞�$C���{UW�.�ոPx���E6F!�z��\���R#4���r��	a�H'�Q�#ɣ,의����
�/ܱGdO����������4���L�@c��&�/[&�=̝)�'r,�Ԓ���������q�.(w��0�]P����ӈR��-�w��y�BTP���4�+���E�l� �G:��R�Mw%�oݗy��aA�#�Z	���:
.ckPf.#?�:�4��ݷ��|����{?���g��_����v�Uh�f��2�<�k����02?��	��0���+����y�m�=N�b�P���Y���i<)Zk8Dx��b���o�6�OO1}�p�XƬ���7�e�@�%�9���X2��Fy}q����#�K_��v�=��5׷� ~���U�����gO4-�r��>�H�>2�.\�h��g~J3��� ����S�L����>8*4z�3��嵷L��A�tbn?�F�۳�D����� �vd��4s�|�SʛtuX>9*��|��5Aw�*�D)Zy&!q�X��ibwS���{9x#1E3b��������Ɩ����Y%'E_*7��f>Q�1�6� ਔk<j�n��d������/p# j�)<��|�Wj�yc��p��>�9�Y�/�%?�.��	��������q�͞[�Ĭ��7��^-�=&ȸ@��[��[��C��X�uM
��4X���&6����g���~~����Dc+��Tx�zY*����k1.�#Z�4\����W�H'44[�_^g�6[9�����!Q_�Mhu����"b���k�0��<u��	
B�#�B��Cݗ�:��/$�@��Jh��x4�I%��o���}tS�Gx��!��S��������:ߕ"Y��ڃ9)�_��>�$2ѱ���l1^�66�^!�-����K�ϫ������
��.-r^�EO���1ǈ|��H迖�Ȃ8s������2�ϒ�
�4k����*|Vτ�+�	R{�UP9����N�~E�{�jo'���K9�蜶nD��^�R�5։7�{T)�w�üʤ2h�p#�o����3	ப�����!�|�.F�U	�hd�N9s;�v��s�e������d�.�8���+_f��r�5�Z� ?��	����u^:�[v�ޙ6�=Ĉm�_�j �-���Y�n���Lʂ��P�����,-�.��U��������9���(u�+�����S�E��W&��߼Z�"�X�핃w0�e�qI���)a�Ѧ������CL�I�����HΒ)"b�fUb�Y��׉#H��i)���v%�q��w�u^��Sݪ+����k��o�s�/�q@�I�ִ��ꧧ�7���i�_��JS�\���~�H-�6�d�0=�a���/5�W���:*Yn�����j��iq��S{�_i}������i$ ���R��1�����۞&�o�h_�R��1P�ha�(<W�)M�h2��� >�u��mK6[� 8���D�����Ӛi�`���mb>ա��&��[�뮢i�ǢP����CA0��l:ر*��n\GP	-����Y�|e�XZ<x\�߷�b[9�Ȅ�¯\��&��S`-�_����Dkd�l���P�&sD�oV�73+�G���߈�7x����B_�!�%Z`�e$&��T�%����V�#
F��6����e"�+e�Wt!(�Whφz��� xaU_�>qF��0
����@���0�OS[�g����d4o��]ۼH�K��C�"�q;��a�tSN�\Ǯ纱%(�<9��I�9{����6Fo��vӝ.�ƫ�1��l����$��=*��yZR��B;�� W��m��Ľx��5���`����{�J��k������1(@�*�ӡ̔C:�N�x@H�\vS�gs,;Q"�DRu���Vi�#��O�xJY�x�8�4�~���.��Z�Շ��҇U�H@e�ާ�
@5��a��U�,M
1T��R�F�%ٕR-k\T�t��v�-6=EX�]��Y��f�kG���)'N�v�">�U�$}q&{�^�Uڧ����'RG�Ԋ����la�̧B-��R��K�G �>t�(3�M�ZT����bV�8��O�C|�/�~�cRCo�CE)����H5s��FS2�۽�+
�Eq�r�#�S�ZoVb�Ь�����)^g�Z7��t/`n�2g�l�ײ����\�	S�� ư355,;��*!��Ą|��I� y�jHc��,~~f]���NJ�\��ј"��]XƮ4�-�(�Epa��C]�7��!�(��?G ��ᕖ��<�MZneD�Ɓ�c�N�/�P��rH߄��NR��Z4t۰O�xQ�i�ӄ�^�����{jK�qK��i��g���gC��6SOes�<2�ߟ�a���<�o��:(,���ڱ0���R�����&�x�_]��H�(0�:�La8i�t1-/y���?��؜z�w�+��.~��B�2>�)��S��:/c�=��C�+�@��Eoh0��#��C��OIȿ��B�A������R�a���$�wЀv��fn@Dۺ���#b�O�N�;���hI�^G�g��pY����eR�p�׀ϙ��G�.���>�������QN���LU��"��,LĹ��lx�s;>�+k�Ň���Qe����($��7:Mɸ]�Oc�ˊE|o2�B։V[n�Y��q7�!��y�x҅[����k�qxŞ*K���Ӱd�_�S��vѢ�>Zj��0��|�s�Q�@��d���{�3��4�'a1OF=��j�2 �����|1Х�N���ׅ�����8�5��A���doa�
�5��ho\��S�G�Y�i�$0��Y��lYH:�3y������"<T�����s��ݍ�B�?�؉���6#ٓ�UF_�]E��;��t
�^�0ƒ��uu��O�s��8��]s� s����eRIB��Ź�?i��ڮ]1-������JPy���JM5Q2;m����"9f H�}������d�P��+벥�`�߫)KO(�q�Z�y	!��d2�񐅝�q������1/R]>0-�L�A$�v���^n!l��3fҖ��]�F�U(�A\O��>Q�Q�Ώ��i���c�xj23�>�w=�� ,#ڭɶ��B -
�8��7n2]^m|��A���LK����� S�mG�<@�@lWؿ�f[d���bh#A�]���ᨚ����ړJ�=����`�I�1�a���:7dN�� ���#Pr]��4��5*Z�]�����u�ް������I�	��PJ�3c����hg��IL�
졔 ���P���+�E�oQq�0��n�n\c�ޅr�0ɤ����@^���xm�>Cч	����0N�<qc�Zr�J\g��a�qE`K�̂3�,�
D4Nx��i�C�e~Vz+�^�3[
/`K �m����,2�z�"�*{XAK�eз�T`D!H�e�}�%he@�O��+蔰*Z52W}S����������+e����	h�[���@�Hkx����7���H��Z>���InE!դ{�]��7��c`�|A[
MwJ��DƯ��|݄k��::���5"<Y��5�5X�T>����Y�/c]Z�<�����2^О��� �U�l!��ʊ4i>�� ^�&��M��6æų��VW�8N/�Qs��o��v%�:�%Ϻ�f�/�jMS��Õ#	�����=�a�2X!��̀ة�IC(�^ԼĢ���`�j�b"��<.f/sn(R��5{�& �c��h�.�i|y���t�� �3�e!T��>HHY�����Oa4�:~�]�=�N���%���n��
��>f$B��:�!z6��� N�$�-Dt4��u l�Yr����P��Y�!��B�<^c�U5$�`�k�h]C.^y7U�>cmE쯤cfJ@���Q�|�o���(���z��Ճ�my�b�,��G����HXUQ�*�Ӹ^T�i;���;t�`R��$���� ����jƠs�>�`9"�l6hmFn���8�������;I��4.��o�r��;���0�dS�x��0�<���H�Leqq�c���i ��x�t��R�0r�-�����g��'��/�nҤ�_���j����^��,,��B���v��@Wo��?��r�Ǉ~�~�*��� �.��h��_���z޶9���T���,�'���r�w�|ľ���e�@䮨6
4:{M�oxQ+ހ���0���lk}t��Q\M�xP��(#+;��"���$h�|�Nϰ�,�fvE�>(�1;��X��S�RT򧅣]��1adR��f�~�)]:ڏ�>��H���.�s�p���ƃՆ�:�㬬rD&�w�1(���,WE+J�CO�.o������Le	&�'=HŶ<�3�I*U�̧}	k��|�~hx��={R,��t�B9���ۄsb�L���7�^iq��"�����/�Ɯ�]��zn缒^\=Q���CcRv����@�▥9�o\�E�����n�b��D@l��>���N����B����"ݳ0�5��t�?ġǓ��S9�� ��E�������z�\���Aj��(�
Ik6�G9tmIaYL�n3��IMb��#���"w��(���`C�ra����{�VB j�x;y|p}m��n� +����(eB��%�Y׫�mr�z��1W	��X�ǭ�	��T�MX�}�՛��&��L/j���_��m��Sl&���E�����܎��c-�f��M�;�-o������[y���z짡��9���/�!���u9��~_a�܅ܝg	T6ڦ�4Lk�9�oN.��8��Tl�H}��D�6ԅm�{#~k��J�k��ء�!��t�9y�Ш٘�d��� �
���Q`l�����qt�V#]�F ����RAJ	�jD0�������k٘�.x�c",DE�'�D�P�Q
�7��;6Nـ�r�$"?J%�략�����'C���Q.���5���_��� IEN.�?t库+��7JA��4�H��I`
����@(�6#����C���v
���W��#�K�:���ĝ��!�X����m�.�9�t��D����_>:�����m���G����V�t�GJ'B�̑�d}�ă����-M�,ƛe�V�L��^�Ѯ @�j�aeP73W:-���_~B'��3�]A.�WD^�#8x j���w��Z�Bft����,����[izu�e�|���+�[���x���^dY�4���
�w��Lo�>�&3Or;1��8�q7��M�ӄ%�`���r�
�ށ��P�t��K�,ld6l,��h=����"�p�K�xF_�yL�Y���oV)�Z-��U����+����ҋҜ�s#�V���ؐ�����ʁ_k�.��� f�����6���g�eh@�*���n��X�>"�(���^��ftV��_ʀ3���Y<7��f۽8��P?��*����I6�q*���n# +�1w�$��M'���i&*�DnL`�����
3����0K�WeWAʺ����,C� y���z�S��g���殈m�����Qu6��=���%�P�����%���)�C4+uR��Qr��Vꥡ2�W�$��g��B�]�6��r�>�3Ŗ�Ziq��'�:lN�!��Hܙ�4c6�eE� I\�}��ʕ�S���w;��Ge�M�\�o�\
K����j��N�k)�.R��,����K��R�J��u�0�jĎad�m�R����TSh�ZM��P
�-�V���N=�j��SJ���i�Td����SzEČ@�嘶��U��a�	�!-�EE����V��8�� �E��8�-D���,���͟�t���;�TŘѯ����Xs��9�(�0M�X�0������ި��D��ԓ� !�xsU�@˷����N��@cK뢞g��X[���%�" @��{:F\�{�E;L�R*ҩw�麛ŗ�sY������ c�����˹֒�R7�	�y���E-g�2Q��iAu�#�-S�{���\��s���!�+�ɧ���S���j{����k�	�M��'�}���D�8�k��*>-��D���u��]��m������T������t���[�s�(�� ���~a��5&��5>̫��
B�����rC�zX�&Gf*���Ϥ�q�6�È��C��'4�¬���㿡P~��1D�ݮ5���Ї�{�T��y�X}�Iw�(.j�fz�W��E[R��.j�D�!�s�,�A�
=v8�S�_%��8��6�q�n9��M�]kA����
$�A�GȞ�Y��q#kE���������R���q��	��ڼ�l����t��1MFW!Y1�K��w�H�D���Ǯ	��s�94 �+� "�q��q"!����)�g���/ӡ�evk�G{T1�*:z�Y#呬�`�w�3��	�����:6t��a&W���5�.�xv����M}��t��#�5�-Ԟ|���e��{���-�+���������#N`�F<��!�?�����yfš; ���g{�Ŭ����*Tk@�0����ɏָ�nv8��N�u`���	Zu�a.�֫�#�J��)�ĸ����H�aP,�����ކ��L��s��yi�0#�Sjد��)���	B��8����T�ʸ����~c��{>-xԸtU�/�В�b��X���<H��n�Z>��0��a�i��4�S���Q���&�q�2��(�O����:f{�q�z_�;輸Q��R?���j��@z3A���8YĈ���Q�m�j��G.3{��<�����YB��&O)N}�'H������7�U��͜ �`�&(�'<�W�����}���'i=�4��,�%i/��$����@�K�����6��sl%A��W��I��0����a-��>��h�� i��)��yA�/c���I�$B�J���������ң�F��q���w��C�n7X�~ˢqq�+�>� �Ev�i����J#Q�wI�U)M��ύq�td%�=��ǜp�c)H�e�$K(�"���&m��O�`N���v���%�;jz�FRS�F�f���g�\�_5���Da��B�8(@�H։#]ͼMa�0y1�a�4�j�<�D�T\(|<m���ؤv �����Ӳ
���>�� q���<�M�&.�KTʡ:e=?�6V�L�:ś�3�
ۇ3���_�A=��M Ѕ�/}Th%08�(���/5��ْ
_a�����@�I��� �J��X�>��y��Yc	�hz
���/0��㹃?���H�����R�=6K�$o"!\���	�=��Ǳ��N����oiIe5��c�f�H�	�YLd�[Z���U�>���#���]��~�Q��>0����6m�fjv{>�b��F�k-��=k�s�|��?r�k��$*���j�0d�|���W+|�O����6}Ř���[D8��)���߁���i���mN��p�1C�������-+FChe�3��#���,#�[��?����l�A4���zt��N�Fl�~�G����Pdu�8©�O[ӏFA0����z
�O�M<a��Mg��1:n9�x�4�wIY�3\C[37�ɴ>�Ĩ#���k�1�Lѷ{��p��PV4����P�w� ��[P�\�Vt�KF��Z~8���+��b��: "�khҋ�N����v��ߺ�u��W��Qa�W��J��bRf"�	|��g��6DS���u�f��˓�`�ڟ�/�������lE���gό��=:����(��G�	�7(�H�XuP���)����y3LcQ%�y©(���4%˲�}`���QY��X\O�L�E"�/T������bJH4X �i]����z�(f����� Y;GS�^��+�H��|9�;X���0���	�������_��˹��+��Eلɻw߱���14*+��G?z�����y��'��:�)?tg=2��~Ss�Xi�"!�<� RS�g���Z�曪�a�T��R:Lv��\Zt��l+(�1(yp�5.�M�+�Z��U�لu�ӳ���w�ar�2���䖵4���Qw�� ۾cxS�@�j�������q���)0G;�0���~o<�� $��	 -D{��EX�i�D��89 ��kDND7�A&Ue�._�M#�Y� dXAv7i�~����S�s��w��|>RQo�F�A��Cl��q��uO${ ����b��4\�|��)��Ô����Z���ʬ��/$jg�0�;�B_��^�2n�M�k���!��Z���:����DC��wJK���o�c_�H˹�O�}U]�����ɷ��n��*�`����+�hkh)l�����v�����؋JKSD�U��g�ҵM��U%�C.l�>����]Dgn
,����W�4L}��F�>T�I�����
����	�4f���&!���mi�w���%��֩�27���dTU@��"#��Ỿ�B��Y�'���"�R)ZI�{E������m�l8*KF��jF�����ҫoJ�%S���,��9ݟ��IG�y��PdM� ~�Q�/d��)�v�A�;->
3�!+�0�7�F>b@A���}�ϋ9��g�"�$�U����u韃J8($���*�����l��q7�h� [��z0ӆ;�<����3�O�x�Buf��@�܋�}���c�h�m2A���ɕjt�xJCsLy��oYx��rܨ����ۆP�ea�Y�1J	�%���Ҍ������8WT�K|*�`4�n�`�Y ��3	W�5�$gx�э�����Z��nY1Vz3 ��;�>t���0��:�;�������
��.9Q	F�����Aw������"�W��3e5VȜl}d-�V�Ы�{J'dK�%�J?��dʊ5f�9� ��ݙϛz����y�`:��Q2"���졛������V�&����E_��1Q�s6j�mr����O��ª�q�>��?=��h�Jj����祀��c�Q��8>���~~m��b�F~n���5���k�=���C��I�{����� UN
(E�}rF<��7�v a[�Sg�����������W�����00/����U�5�)�6�����!����OE$2������\�R�G½�Sƺ#�N�~n��ж1ökQ�Kr>��l�<n�h�*�c( ���ۊ�0��Z�(���vM����A�N&�^;I���x�-�iGv�#둎9���H�����}��:>a�0T�� �f���{�x_.�Y8�
̴���f٪H�Z��T[ZE���H�lJ|��K�' �XpKC��"VW E��%V$��Fm��f�^V�Q��*�/�b;T'N��{�oWrz +� Ża/A��a�v���""C?�,Bwk�N�2����pso��-�2>������2�G�z2�^1���%�:r��!*su��i*Q��T��,(�1%J8F��B�3nN|ܝz6 ���m����2J:QZ`e�U^	o����7&@*cm���c޲��Y�'4H�㈞�z�\KЂ�b<�&�'�w��mظu	�@��?;���[�����i��.�ͺ�Z�|�5>�E,���1E��+[
�2-�2�rg�,�4�5Nh���1Ǹv�����n�����`���#��}=�[�#u��A����`���;��{������b$$=�1��7m��S��<��L�s�̊+f��6 &�����!�#��K^��yt�<��`��a���'���'�D����lގ�p�p���L�z�JU�E3*n���vG�q���O�z�t�%��4�����n��S�q�G�G� � �hw8�3��i*��_��;���S�)l�^�;+� ����n?��y{sP�E'����r��%�iW��6�=3���$�1�}wH�H�G�QVai�~A����g��AB㖣,��u׃�R�N���w�e�7'��7���U����6�{�Q%�{��R��Eg_
�)��x�~�Ȁ��j���',�n�H����2�O(��4�d��9U�ldU{�ӄ��D\�E���")���&ֲ�w��	�*;\��q_�f��-]Xo^B.���i�5���g�Q]�;�%�;�"YNmT{77��n�.�c���ע�Щ��T|�[+Ա5(uV��!^���)-�j��w�9��%�9E/�q>?��$�|��K��_�� �k����W�6{�LV1�|�)��tj���K�ن��v{�"�:�ؿq��$aQ�qP�\)���R��gX�a�����5`���$U4r�&��Ƶ_[������ٓ#��\j����O�N�ϡ�k
{�+%n��]4i�RT�7?��O&.�.A�(
`TT ��kk]F�=&�2�s�鶎ؔ�@kx/�+K�W�,���id0�P��=��e�8ǋ��UF?�[�'NiP܀�>�`;G����r��Ǡ���/.��%�����I��Y$P��ٝ\� {Ԥ/<8��?�I��;�!h�����-N��0��s����lq1;�̈h�	�i~=Qo��Q�~#�&��Ck��U�M�SP���2r�A��y�,�Y�~ōh������!%�D�:����y�)�"����:�(�����9��L�
6۰�?�Y��]��0f�q@�g�K1�v�A~	�Y��u, k*��f���8k}Zuki��D aӘcM�f�1�pB$�ux�kO�璘7 ��!�Y�ۭ?�7w��ō̟�@�vF�K��� ��m��{�+�5��3��ȹ�t6%)WG&F[j�>��]�n"}���R��e�M{��}.�Yz��Ģk��N�Q|�&̛'G
�k]C�,P
�/���d�����IH6�w����7|�|2��9	4q�S7𪂵SX���,0�̧�TZ��8��E����!�Ds���q��	Mq̬��W�uX9@��&��E�x ���+�MoIgCC��b򖡪�yl���t&{�'}�1E��^q�0*�ǇmU6q�PA��j,��o��I��DL[�T$�����i�]�!`��p�t�2U�ec��'�z��ʳ�'���OQ��lp�F�n� �*W���HJf-J��f	;�z5&Ԛ#���$�����.���1��m5���㹴E9��R��&��#�^ά�6|2�$�QGA�p5u��:~��r��)��E�XO�����>n�f���ީ�QN�ӑr�$�1����-� ���:G��X���ɠA |��
d�����s7�|�M��}Pdd�24SR�Ý�Y�s�!W33�,U%�g\ �A��L̓P������V��C=�#<e�6T˘X��{cTD���P����3�1����*�7� ���(�S<�p�=�Z��q^��p���O��zpu�2k�Tԧdf�W��Oʶ�>�x~`�wm����V�D\t>�CŔ�U���l���?\7�+~\}뇃%]2�xWy����/�Ч�ek3тE�V��Rh�4>xq�e��@��Ed�
��B������:�jy&�:�=W5�h�p�0�Q��jF���?�ey��)c`֚;!Lj(��hLrh�ɌʞS��|�$�vO���yͩf	�����6�C�Os�͚*�o���a?W��Y%cM�h���7�!+Hb���BP���ɂ�V���_r6�D�� �i�Ri�{DBU<�\��XD�xz,��g��ó�Wӆ3��cvG���ʊS��/K1Yd{��������ˢ�u��ԎW��X�4�����jjj P�*�x;M���x�MIym9�{�����=��7����V�L<��:I7�� `���ѫu�C"�m'Q��-��_�p��35^��r�ӊ�m 7�z�
'��5�DL �)mш)O��F�k�	��񔰨fT6��A����J��x���v�1�ao���+��t:���a/�w}FT7>0��t�;UJ�o�V�q����LG��%{w9v s8h�#�{i_�J������Go���a�8�T���{�ʨCLn��ʫ��" DЏ��cL_��q���m��R����G+�on�Q��Y�2QeC�Z�(~��dw��`�AZ(�뚤h��ٗ��ZbK�F�y�ns�]ċ.�>�m���+vd�� ��S_P���֎�O�qeǢ�bx��7ԗ��?v����@�ې�-��;6DK��#���c�i�nR��IHG�K��Xuu|��>����%�~�q���{���4:-���,J���nԏu��:���U<:���GSv1ha�W��g�nƠ�H�i)Vs���lQ[8&2>�N��!-U�.s���PK�p�fwaX���5�����H`)abe��1����}����r��u�`��_�%�N>�&L߯���AW�W�r�XY8�!.���Xt��B6������C}ĝ� Էe�Rcmb�<Νx��K��0�{��:C���JZ�äuJ�w����mدF�?}x;EP��!euȯv-�_��k)#�W�FW�rS�qyB}ͬ]H6�_C�
�]�8'C�0�Ø���^C��)���C���<���3�ߟ�Z��+.M��%[qC�X�XZ�*�=%��(C��h�� ��"X��`���'��x)ѥ|$\gcQ�HB����&��]Eٕ"�@e�C��:���wpq�4-(9ꬷ��R��%Ȩ��ː�U�!�~�P�v���Mʛ�ݩ2��dL;�Byl�>_9�ij^�npk9	�+;���J?�B�m�'�7ގ<�R~�吰)��������}!������#�KV���L�8�k�sY}�m�`|B��f`�d�.6Oj��-z
������:����k�������O͖��L�|:R)f��(�BΖ/<�6p�������0I�_�Q�J�hՒ���un�^��7�����w+�f��`��J5W����ԉp[�'�h�F'����"�ȥ����0��uC�?c|��`���g�kp�NϏ*���p���c1�V-^o�iY@ւ(-�w�k#Ρ�zO�N�H0D��3��ʮ��U�̧G�Q�	n�[A������'RQ��g(a^�� �*���AY�wc�G�._���'?!N�[��� ��W�L�#�0їg�.���;Y�OXɳ�@�u���N�����L� g�.j���%�B��l�w�1��h	�e�Q��3���^�E�r� ̘=,�ք���Y+\��~��r�{�Ơ�^�m���I;��m��B�*Y���욢�M�vЄK��p��<фf�j�|�r~<b�3ۃ��B
�~pcմ~��R��nXF(2��$��>L*۳?$�l>I�N�j2��1<ܒ�)�/�ѕ�D���{����16̓+���]8���2�B;b+R���TvI_�RfG%�"4q
���"��4�\J`ӻ� ��t+x��=����o�	K#Gy�y���ۇ���*�+�lB>�i ���l�tsc�^���3Pv�n��{t�K�s�u�G�h��O���hHL��ә��8rL5/���u@c����7�+��d+��5x�N�+�\}�Ci���J���6�c��?���jzj�0���<�>8!.B~���2զ!DB�]@���b)�%5���0�"��zD/۝�Պÿ�G�����ғ
'��7c�x#~Iʧ{�`�
Va31�Y��,0��C~��;�t�\W�>
o�A!+�F��4���x��"��p��кװq|GFK�g��dd-�r��*�}n^7x�x��N���ta~���Ծ�o�:�TQfǉJ$�
���P�hz�-���~RBW÷��n�5kaAQ]��� �<Y���MW�,�]ZME�Z��'������dg��S�����&���z�W��"��F����U�h���������{��0�{��١z���]x����e�n~����p��w�ޓ��fX�����i]j���Q1?�� 7��NK��lt�S8��݆"� �E:J�t t��ԹH��Ǎo)N�D],]�;®�/�c�z}!3���P|���`��~v��ď@�q"����?��
�`չ'��W?�����,a��1ٸ�&���ӡ;[��qdz܉���u���l��~-Z*��M����B<\!���BL����s	W;bc����r��;1�`�)K�CX홤�R/jE�_�#r���Ǘ�V��i�?Ί\�+�ɻa��2#�~��-���Z!r`����P<�	��/��0Z���&�_2<#s]Ջ���7�c��D�#OG+��?����c�߼�nj�wA�ōU������Rq{X�eN�JPكjԜ��;�����zRc�{�I�!S����I�+b�q��[:����ց8^�ڪC۱=ӗ�=�����+�k��~�Ⱥ8Q����%��η�?Gb�����9��9`͎6J�0-|ߢ��j�ZTJ۸<��a�0�Owt�
��;z����zY�/��R�)Hk��"�>�X�(ڴ�b�)pS�f53��|���	F�xXG��{�/��
L}1�90���~�-X0M�բªc�� ��]��jf�ޢ�o���G��f-� 2�=��=�$7�i��37�ȕ��)�/<5��rS�v7�o�jE\#�S��d��*��[�s��1tʼl����J�,�3"|oy�K#�� ��o�=������ܑ��ތ�A �����iڋL{ԨW�R���Ā���'��}���Q鏽�^<_�q0��oYn8�3�L=H=a�m/+��O2��e����^�p�}��[J��,�*�~�����/��*Hl��p�S�#�rM���o��4��}�ȷ��;��F��w,e�XN]Q9'���Vڎ�#`8(`�.�H�ѧI�����֮��7��*,��5:��Ơ��+�.Y�r�q-խ2D���gd�蕂
�1cl�'���;�sF���q,%���/�ǿ��l�|D���5US�&���f��0�\�ė���>;hIhu�̮냣lS����^��&��Р��Ȼ%Kj.1�r;h��'#��!ӊ�7_�1���jk�����+���d�S�zJ�hv���0Nɇ��E��:���%�.o����L��-�MѠ:�	�è�7g�� tu��	@z�e�s��P��F�� �BX��Z���"�čEg7�s�h��_sI��	��!��.�v����`T����ph�<C����Fr�\��a�<n��8��ȵ��΍t��RU���
�У����ߏhv�_�5;*���8��4��qŚ�oAL�.�H��x%a˪P��k�!����yTV��J�\�%LYW�`�7z��O���Z�#�=�&\�r���eϒ~��yW'�U�#�0i�~AC�m�f�����@P����tO�Ѐ!���{+�AcuY"Z�"~V�nФt|� �c�i3W
��s������5jU�����뱳�������2�0=����]�?��&2fI{��$�?ԧeJ��tX�j�-���5��:)��4^�-}lh}&���[֌0=�q����֞�u�hA�S[f�%�wKx���>�rȨ?�a+y�ޡ�����<������<�cB1<�8j��K��֥�oh/��8܏�{t�-n���I�~
/�>�D���W��N�#��B�h�-o6�}7ʵ�2 �+�7r��w`x��6�ڸg��ucn@2����3A�!řBM?�k�:ʛ #uz��+�JL}D�?��|�����(U�r�/��AZ�L�6����|W��>�r>99��k�%W k����}�h���?bD[9c��ۨjs���*%��D�"�Α	��{�PF�E��ۻ��C�~�Ξ�ۍ�)y��u����K�V�Sg_�]9��^R7N0Pw�mn���V�Y$@��f���AW�1L8d�}_c\"<�J/�I$��F�Y�h���J}�=�����a~�4��;W����	ρ'�ӵ��t%��Ϲ�Y��X���Ӳtd�g �ԝI�9Mj��J���F�0���'�@�eΩ"`��CA�\�^�~E�n���樝�����Μ��[�e�J�Li�\��wl>H�l���my��I��e�(�w�����n|g���j3�"w�K#SL� av�^�}YNuz�h�r)���D��h�O��;b:Gt*f2������jyn�ُ�*鷿c�V�/��'�7�Ai�adA��RP�����)���������7���3�P�uo#c��5����^��:E�ƾ���څ�t,N�u��͌+B\�Ɏ༰(���F��j��)u�Y9����p{��.7g,~ ���$�#�Һ�<�D��c9�����|��m��8�{54/=�C�o0�>�Y�v�I�U�T鐅z���M�� �n��3K�3�`��e�hz}[�VS��6�d�����n�T����qM5ª��o���oE�g�c�10Si�`*���$v
�S7���n!'q�m`���^r�o\�J���Ij�,VзmHqs$֯S�
�I>��w�E��~lp���βp���;*�[�<M�:��(��a�w��hI4��ʲ'�k(}i�u��ʼF��G��Cvޚ�b}���ڃ�K�"��=fF��X�H���:����pZ����O1D����Vx��z������MYY�Bn�lԖ �]+��_@��)
�<�_��v.�m(�"�3��X�����^�t~��PD�^C�m����{ȊQ��!��2���ND
r�SS9 ~��m#�6�xٍ�à�w>Kt�?����c�3��E�g4�t�a.tq����*L�\+�DBQ���xљ|hdg�G�2�kW������oA^�1v�dA�{^\'f|��3�NV9�C.���i�9Z����, ���q'e��\mW�C��\�|Nx.��|�����M��_�5{U�*�J������&���Xe�*Y�� ����3��>��D�dm�*o�Q�l�����"%w<��f���C���=?$��_|~캡�}P5�0��u��#�!���P0��;18�'��/�v�Lhx�*FJqo=�,軓�L��w���>��@-_ho��o3n�*�»h��o6GDԅ�+S;B�
C�І�3g&��U��Α���cF���P؅��oq ���6�[��D%�dŷc�����dx*f1�d2bW~�&�8y�t�K��t�Sg0<3��|3RA�<��XKƮ����
�_ޭ�/���҇�W����+����lf�!w>]�G�G�Q��ǲy����:l�!��܊�-1:�An��5�J�r�:��%Xv<�D��M#�+s�|�m�ŭ�d�z-��ai�����:��ŧiT�{��m��U+�uU�[�E�5��F�}��{F��m;�_?��&F�QK�1�rT�Y�a�aTjR%��nAY���0ݍϒ]�k��82�$_]E�b���gi�C�i�����w%�.c�D�r>�QcW$����"���j���M�g�xz���B���Am���R�El .��I�ċ��:����[��I��ʤ{ьcAmh��%x�W�Z��t:0x�o�:.�p%�y�[�~���?�/ƫF%[e���k8�,�d/F�h���1l���c���������%pO�����g+�U$�ڜ�q��]�+�p��P;�$&�9[��r�ֿ9"�ɷ?a��V\�µ��0'Ҫ�B|�>�b?o�,3ޓ��B�A�E2���fN�i(x�1����K�,�J}�B��nbr<�n���|:����O����;��ve�#Co�
���3L�^�k��Y3N���n��Յ��l����� 1�.��A^&�WL������Z��x��2��g����wg�(�&�F��ݗ�Q���g�p���`�;J�:ٞ��)�^�x��_�z��tI���<�θަ����[�s7���T7�$�C����m�	珸5�F� �W�V�R�7�W��I�9��Wa���[O� S� �.�W/uw�Z{�(�HR|�t-�'�k�_�۔���I׽��"��D�Ѿۉ=K��*!��
Ӫa�)��|;� ��L�q�9�]��c���\�<�!#jSx��0+��ؼ�����hF\-��CQt�g�M���t��ƚڎ��^1ɚ�B0�Evq����Z�����$�n.�v"�B.U9K�%#ҋE��	x��1��E�����k_��cq#~dГl���A�ݧ��IجB�v�'a����w|�����3z��^�$g��is��$$���iY��7EJ��s'n��� e~�i�7Bu�t��,��+M�%)��k�հ)�^��ozZ-��,ꘇ�ǃ�j�OA���ΖG�+�j�T1}�<?��n}��8U'ћ7e�۾�$J��8�Q�Ԧ$s��߲���?M3��@ِ+Q�����?�k�#\1%���-)_���wF��@m	�e�o2�s���=~�z@ٖó���(Y�D����mTu���� ��z�TMu���q����9����۶0��C��|�E����\�/��;�4T�*�b�
5#���7-<��|j�D��U�y�41�h�C�c��}��W_���hb���u��0�|W���dK��v�]5C�"�R�f2�#�q��ڔ�/�LS���ώ��p[�_e5
���F�V�7�J��"�/hV��E�>�ǡ�	���P-]�z�c>3�>��iB+��۪�h��x�j�퍪Nk���S���9ӫS"���~P�_!�J�S��F5�M���ZN�O#�F��Qt&��$*{pOQ�>���� yՆ+��7�uO�Qy#A�</9IR�Rw@���Z��9�Z�� �Z�;<��#lΊP�iJԮt�H��T6�T¾h�}-a�5\���
W�ҽ�	�'�%�T��<}�ʀ�yMI�{D�7S�+i�ݟ�<6�M���>�FZ��ɻ�_k�6�����b���K<gUI�V,?�^�m����1�5
�B����x�Z?�����H�P��@�^��A��l���.c����'y�:��u\�%*��r��A~*`H�F�7�7Wү����O��MF}�%�u�%P�U��H:E� �L��2�bI˦�'Z�/:Pʹ��+lZ�~�m�K����>�\�An�'�����I����o�$�����a�@�}�Ԋ�rw�g&<Nw4��1���zZ�(4;�^��������Z�n��m�PXF�KŌ�<�v���~�['@ٚy7���� L�	6�T#>�}R�+���*����<����qPK����Mk��?�a�Jm�z�Q�������`���@*r1�����bZNU����1]W���C.,-�%&�'�s)�|h<�O�4U��$���7�_����j�|��+}�l-v�9�F;�,_�vjELF���ɱ�2�k�q�{��-�ݪ1��R��F!��' 9��b&=�g!��}OB���7��k����rc��l��vz�'4���WM&{Pg�^`v�����2Nu��i��2l���-��V����h���@�W����t)ٶ����5Վ+�>(����y�
C�,w��I�5�B�h�±�Dd��
@�ц�*�Ki#(��&}��9��u`���$��R�����m��ta�6�:{�f�R�qT}�^�X��� �q滉�	H��j���;�E��m��+d���l0�����'�%zU#aL�%�Zř��������svƳN�h~\�w+Ss���H�_x����;yb0�K�ƭ��fC���ǈ竻TP��ks��&�W�ڔ6ؿAo�zH���^��F��jRwUT
X��4���Շv�Q�{���K����'{ w#��k�$	�1ΰcU9�,{�H��ރ$�6o\9_O��/;�K��1��Z��O�u��	E�0��)�wD�@���N�|�+��Ox`'���c��BFU���W~�_"�^T^ρ����d�#�9����Ej����$���nǘ���|�Ym���>����%\�h���@��;�11q�6�ų4��:�t��_Ky6��?�(!je�
�G��G�9 ���c� �)�Dh
��s� �aK>0�	�IO�8�Ԍ��s
�� h�S��p/>�&X���h-.\�>��?��T�+1����\9���%��ON)�>��
��ūf���XY��*˱/�6.���k�	�}����M�u���ؚ�'s] %eק^l��&PLށ�ʑ:V5[��"�f!^�*K�{�G�2g;9;��Α�����>q\Y���c�� M �-ea!���o�::U���T��I(ԆE�y0VRPY�_@�y�F[�(9P�������T��_�[������O��|\/O.�U�Ǳ�
(�j��X�3i�:����f�^	J����%�X�7��S��[#���hD�{q|Oɡ����̪��4�+j�^�P��Bh�5�/]����U�3|B�89{�gr�%�3��@��8�Csa����i�gʗ�o&�Dh��s�&��_[5�=;��|N�7�\��Cxa75���^��OdDl9�~W��:	��RX���8l�~U�>��Zêz�� ���*g�ؖ��?�uM��L������<�{,�_��Ӯ��k'B֖�I�:v+�x��'+��ܸ�#�YyZ�gl;��y]���-A����Z�������`#e�M~�� K�u�&�Cd2�w2 d��k����Y<�^fO3��EwU:��7@.�/� W�Z�D�-1�-��%hə�hQa�s�6A�t	������n,n(�h@[���/tt�12�z��wA�M�3�.:CmE�
N��֧��L�hJy�AmΡ�Ʈ$��j�4iA\ֲ�Z a�~�Vw���"ڟ�XE��b94P����[lǫi�+�_}��#ר���� Na^q����K뚅�d3y4��+��$�m:�r�=n7�x������3�+�&��]q�R�jAR�pf�]H� �p�?S�����u�5mƕZ���y��F�Jq�����Z\�O Zh�� s-��/HV������`d[��I�y;hEloCǹ�&��n�Q�1��O�8N�[��
��Z:8�D�8T��|��b&$����z̺)`�|�_�)g�P|��u$d�5�mK���Y�X�����Þ�$��MA�6Ku)b��A�fJ��Q�;�mQ��'�B��+^���v�~�[�Qݔ�7���jl&tv��".1�\6�]<@���1GG�{
�di�@�$d�-SWn(#�j2�ش<��iG�$ֺ�泩\�`�X��Ψ_ޡt&���a(���z@�hϸ�?��
���Lp�kK)�4ǵ���Lᰫ'��-lw2�e��p�ٴK���@>�;(l��[3h�6{�O.�P�	�6JɈYb�eXp|96x��U��7���_Ww\�}O�!
�h7:�W� �>�M62?��T�|&���a��!Sy;FBA�K7(�kj(z,���:j��WpfI�xe�/�}��$�f��k�eU�*���<;���x��I�@_O�8�Ձv+7QȊ���Up{�ѮC�L�n�{�S�J�k���R��r��,٬f���a?ė�dS�٤�f8�*��gU[�1���$��/�d���kr��̜�_ɾBų�-�<@�oUM�c���J�H�[�H	]vW����	dnW������Ǔx�����,��0\7ݶ�X�T����o�+��s��Bt�!i�����ds��<`n���,)� �Y6���ꈑ�n��S\������r^�U4�Cǆd��2H�i�~���i3�-���M﹬Ģa��@�(�c%���(�V����&�,{�D85��kF�*�J@���x�G5K)
���^S�v�`�8T���T�'�3��+�y����ȝ����ʣ��$\��6`S���<�N@�
b�ii��&�)G2u�/&ύI����TL�������p0��IRX�E��}ET�*�یF_@~��ᦵ��MH��168�#-��mE������_ݞDYK���4������#�"���" �f!Ꮀ'�Hq�u���ܷ�A�p�=ASN�f��/*?� ��\@坑��yn�����d�!GͥDn����ÿ�܈\�E�E��w��������H�Pw�3�ph�]�$T?�y�}M��c�#����6�0��mЈ�:�����Ao�b�D�����Q�f��z����d%�b:�;��H�2�䇦qN+�j^�8�Yy�y��ڎ7�.�W���r��v{��@�B�Qyl�ź=��"rr���Z�7������K��D��k�(A
9�2u���Q�Hj>1�;����	y�PKj˷� �ol�=�kP�9^�2��
ny��&���=�-����L5�(��g��i�®���8�
KE=D�="8��Du�Z��*�l�^�=�d�D�����R�����f���%$)�-wl`��GP��nwW��}�/P�eX����ض~�n�`Ī�_l����>���9C��z�xZ%�;��(���X�˾5���w;���t�@�-�%�ؐâ.�ue�N9�J�"zΑ>T�t�(���9�C?�h�n�]�Ak�Su!�����/��Ϻ�s����mu��z�jbs�o���Z�8"�uT$����G:zi(�*�~9���+3b�Y�7Yv��c���|�-�R��f�|S�<8@U۟�k��5�!(q4�mB�9�.��#��s ��"����18�R�^j����uw=J���^xJ�Yn2
B�!�����)�J������q��I�E6�V|���[�)O'���Ͷ�����b��o���_H�����)�{��p�Xq�Ĝ6�ot6�5"{���]ȱ�K�-@��,��7QӉ��"��q��)��s�(��ν`uT�s��X��4
���[A�%�2xC�k�8R��� ���䵊;�x�l��ʞ!���Bj�����$@�4���	�$6[$�A�3+�p�� �}��=�:BL����C�o��K�+������r}
�&�uvF���GV�=5 |�߯c(�5 @%�^�}1�~L��V���n�y|�Qkͣ���6 ���w|�����Ym-���fN;n%v�>Y�a������is�1�KMZg�01sX�Wdi~J�����I�mce ���.0�M��X��d��f�zu��PyC�f�YM��[U��4ۘ��ni�׏�m�M��%���p&A:��#��gw�b��k�QN)�bܳ�`kTX�E��A�ɉ��Ǳt���`)���_��B����%�I욖?����&�b�3�-�
������0ri�|�"���}v��W��!-:��\|���?����W,@ ~}r��EӞ��Ղ�T�跾=��t@��X:6d�ﱛ�$�5�|e���b�Iw[�1��&}�6���|�u?�&U�����,UV�mQy� �d����]��Tb8���\@�Q��,�_�_�ob&1���~��L���9od؂*gA!P1�#�G��q�>e�WI��O&�ǎ%�V�]2�T����M�QK�����^Эs�������4���e�jH�;{�fl �� ��̉m�)����3giKsҽ��~w0��%��F>B��@���$��ơ~Sg0���X��+�}��Hy��9>3J�
�b
Á,�vm��@,�|������!I�g��B�亠�)��% �;��	<�[N ��fS�פ���1�ô�7�ڪ8����Y�����j��6�_яGSM�v��:{�2��vea*�Ǉ�9�}��x:�����i����?@�	�cM��	¶h ��:��Z���ۨ�Wd����59&J�Y��E�8�����i
8d
�n����� j�U����R�#��������H.U�ʷ�=�5���2҈/L{�PL R�r݃���@xM�$88��)���H�}�j.�]��V���m2���(�������Iz)�OJ��������/�T!��?λ�"qG�^�lFn?	��c�S��̿N�kiƋm�B9ۯof?b�@Ʊ]}V)�c ��0�K��UR1>l��U����2�^�y���6�g6�@g�q�~7"��������L�'�_��vbR/��O��yE$�6'��~&��їꅅl%�f��mn珮ka?��~c��6�u��z����@L.a�������Tr��f|��Gt6Ѣ���?����}E�K������q�$)���D�F'4:���CĐx� ������������#:Q�v���l�2b��a�������^˖?��C��~��Ɔ�Q��]����$�Œx��ٖ+�?��f���UV��r��l��WԨ�m��Aze�ROP��K�`��b%r�������)π�lZ��C3]r�OL��f�.��8j5�$��m�A7�s�h#��%��1c�傴�vԧ�k��N�M�5e�XY�dQG/�����{�1��$���7o�g��yOwO�*�@T���pJ�a&_����:�*�w�ՓLD��xg�uy/�� ���V���?7Y�"U��9f��e����Ra�Z�r��C+�#dhNb̦�*r��Tr�.��Uo����y_���/���<Bz�C��󜴈��n�3�Y��^�s���*��q�eB!�]C+�VJ�n�y��z��k�� &Ɛ�P
�;lg�	0�����|��F�jG���n9��CX5N,���7�~rq
nN -=���T��������	l/���c��QW4�im_e�۪G��_>�J���m���C���Ua�Z�M(p��9�J�4=���%q���뤻'�D�sIS��AUޔ�&����F�AOʬ�2Ԁ]{JY��X������t"\q��q��h�yA
?���	����(�C��Z����d�����}G&(m�ԡn�� ��*�(�*��^���m���]�vϱ&[t���`��ߥ����Z���e�h��֫O�#���/AF�\E�d�v��y+�rD�UgL���@��g	��':�<��$�>��ژZ�Hę_|}v����&���\������uH��s�|���ԝ:r�vo��l�e�8����@���jh4�լ����H;f��V�{�od�iI����U��\��2���I���m�

.{����X8a˩O,�����SiO+��S��ԅ6��z� rO�]�P9tF�˒TDs�ƚ�H�u�p?�I*c��$h�D-GM�F���x3�%º��W�&sH��S�kc[7@[�i�r14��3����FC,	�3
WAB�9��ahd	��]Dr��3���c�k�* �F�c#ڳ�"t�w7������eVj;#��}OW��Ȯ�
a��e`���f�Ʉ2��y����t83�ru	���ˁ]�ĥx�����*JL� 	���ЂD��
��t��Q�4����V��N��C!X���v����~Q�mZZ��ػV�i����b�a������⣁��QNެ�y�ֲxdޘ�� `,�^>��\?�=�l㷾���h�%�r�>�����*F�U ������	�X��J��6N�Z��֟)7e���ɬ��:�A��ń��|�M�UnW�ţǵ�ІS�5��l�����dw��&��b]���+�����$Į���mn�H(�ޢ�u���f2;�0�غ1�œ��)kZ��aMӿ#����.$�n��~d�	[��E�Q����
�Rƀ[y���^���!�ղqdK4q�Rʨ��Qe������GSv��A��X�u�:��ㆧ�y��~ yt&h�'Y��b�<L~�)9�����M��`c�y�4����=�ix
�����Q�3 ���XI�'�hǪZfͅȆ-�}������Ϻk��UF%9���zbr�}�N�m�K �Rx��Ql$��z���k���=�}�-�.D6T:ɇ���ַ;��z��|St������FJ��w���E�4���3�T90������[K#;�`~Aު[���vz�i����$0���u�7K�2'l��b��T+�����}��|X�z5[m�^��Y.$2O6嚯�S�Tn�'u4f��c���/�ὴ;!Ԛ�c[Lj�_�B���՘���+�w�b%.�~;nL��PY������Xp�B���v2���y����URƠ��4�����M݈�����~هbĎQW$�d��v�X3G�</2I���,s%���wz$�}�}����d�x��䴮�
Ǿ�k�v2Q^W�����y�e�'���;�B��U^���ݬ%�=Ӡΐ��sX!��>��\�	u��� �߼�0�a�D���E���36W�/kӢCa�"`�����-��]r�A����G5!֥
H�+s�9���������2 6��6v��({W����n���6T</O�a��+��h��&%��"Q�I�ws�ܷ��gIU�u��}��觃�S.@>�R�C���3�N�Җ���Ĉ:B9�\hVʮ2��M߈:�+��y�ˇՏ��.�:�}��&1��0�hs9t�v�
F�O�H-!Y�����8)���b��䳥z0���?�T;r�ے,������s���|ʘ>c��6�.�_}�q��ی�-��Б����u}�ȭ9G,KK1�����b%�:&���W��0�(�O֩4:{w Tբ�e��&�QnNy���*(�l��T
�2�s0!���{�L��VH�B�m�L����(>?1����.�M��)�)۠�R�3�4��DrhfCm�]�41�[�}�ם�̓��AB�����N9��J��^-¥ն�y�B�����#ۛƔ%��J�7y�"��.�����ŉBDA�xpK�7]����~�(��[H�[lrgG��L����(��!A�bǀ��\�)��JBqpG�l	�x]G�U5�YYw�`O� �XujE�O�d�_�����d��1�ME�MB���Ɓ����^Sù���t�ϻ|Rd�r������
�����7=�_��B//GӍ�~��`��6�^n��b��T[��ɂ��i�a�ly ಒ�]x���-₡Axъ㕁d>%�f�3���4E�ǞQ�b[�����.:,��^`XR��o��ac�d.\Ǫb=�����D�QTa�^�쿺.ޞ�R�m��XE/)]�3�_����&0�1�D k�]��.�z%T��#~�G�-��$��|U-��H}�ve(H=ZE�+����W2��c[bCG���$F�+��<4�9�]�1�#/��@(�{~b3��Zng��l�0��-��{�g�|�$�)�I�;@�y�7��LM������������ȉ�͛����@{y�� Tޅ��gӦ贶Dw�b���E����$�<��-��qeX@L]���'��+�j���^8\+���}�\��(X�Ag��i
c� ��E�ҋ���d�یowr�	��1G�ф�:D�݋����U�٥�V��5���#�$�hא[�o��K�<<�nO�T4r��,���4�>������9m�g��+K񯬻�Y�'�ػt�Q+#Q����\�Z- �(왴�C�*��m�V�#��{�n@���M���^�wNzdF���o�H��t�-e^IC���?��Z�����ߔ��/�f�x��}� �S�HMET������)ёA�u`t�,u7JH05�9����'�/�Rpo����&^1*8��e�����&��7�ė@�
CD�/
�㈏�)TSo���k<(�T�.y�qU�sIo�.ݮ�zHi�ʺ�A�6�މ`%B�����
�L�Z�����U�䖀����0������\Y�v�.?G����c�ʟ� c���Y_X3�D����wD0��><��-�o�a���Zp3�����ȍ��'�$��/wOe�5��C�.����cΓ�}�,@O�aH�
�Dl�|4��u�LD�=�����,m�R�(�&mtC���@%��v&��U"�w�����c
K������U�`5q���{�B8)�~ ���	e?j�6F֔�~|�,�'�k��(�����1�HDi$a�!ur�#��G�>q��@86ˇ��Y�*COY��ж�SH�����Tߍ�����$C�zr�Ӥ�/J��~=^U�ӧg�nT�c�F<>giF��$�~C#>>����	J
x��<)40��s��w0s�/�@�(�������^��� L{Đ�X��0͕3�?͇��&��-.�fۗ\v���+�[�z�������^����EˣY0��+�)�f1����/�,w��NӾ�rF��؊Ɯ��S5d�.{YP�e��1���5{�g5�?Pl|"�֌���u� �o�P�"�i'����x����J���ɟ.�(�M��3aJ6�M�ɡ/�����ԩ�GP�q+>�}�^�-BՁ���o0��,���+k���2�	[d��;�y�G����I<k�7> �B���c�E췬V����/����u�^I�U"�]JߐF��[�CIs�6�A+�����|7�yB��&�a���\�zE��!�����=R�<\��6!t��T��N� �%>��|QɘLOQ]����QeV�e��'�{�� �s�vВU@oD�X!��<�,�7�������=_�������^X�gy�{k�O�߃~�������l9�bO���SՖ�ћIp�U��a�˂h�E7�%r�K@fpkS��bcRL���I��k��נ���Ҳh5�kl��ӹ�����o	]��:�����d�Н7ǳt{ڵ�@�u��=|G���h��rk���#�e�Uo}1��{	E��{�O���K�b�>�0�:��s��wZAw].�>J�v��Q��;,q�/^J���v[�Q!9;�U����ˉQo,c��m��-�)�0~�.nskE��=�i��I��y>���"9/�E�Uݗ.�I��)��8��pH��,���Ŕo@�{�wVe9kH�ܑ�{i���#=�l�X=�Z�Ɗ��D�雪p�P����"06j��Ά5 .&t�֡g��6�P�N���\P!y��i8q��$�a+��&���ak�N��N�)_���6�sM����mZ\_���se��mu;���u	s1Y��=*���uٺ��J�%�����K,f����
4R7�]x�rA7�c������+N_���ʊ��d��4�.*��S�1b(ˀ%���V�+� ޞ@.I�l����,0S�1�CH9M��E����w�6�����5�{6���؟;ZY��0���3����ӱZ�)N��s�Q�쇻��,�f���-��o���8�u������3���d %�YL���� ���y?�h�P�h?�G,��:N�3�NW��J�xo�
�v�\;��#	�s����1-n#~Z�gi��E/pc��\�������v/���p�	�M��8	|ߟ�V&Ci�<��F?���A29`��+�R�f����h�>��Ҵ7���c����5�a~�>
��~�KPMF�k�*�nЙ�:@���3�g8�-�p�.��Ǔ����9x��kl���b3o/��~F���<u�I2�^��l�r`��x�7���6'=�3巉c���!�-�t u"Z�B�D�*����6�A�&ϔJ�_������U�4Hk�G��qUa�Ϊ���;��T�z��eLr��r���3�����^9��hH�}3��B�kt�"ެWE;��?%dYU�Ԕ$���h�oN�|eI����S2�
!4���M5�
E��eP9�2
��:��Ϗ���-��-~J�R/%�(�㳐�T]����_��+1t���)�RA�q��-r�yx����'k��>n?�sz�SCW\{�i%���X}z���	4N@$�B����[~+:�W���~��$"����sj�>��!$���f�xp�+����y�'_���J��χ�0�ӫ$V�W����%ҌWb�N����7�����sv[i�U�.w�ߖR<o�Y��B��`��N�(	'K�������7�%��Y"]�v���UzYW��[�v��g���7�-���J3כo&;�F��>|����؆g�[sY��̅{�\&Y�^�����02� @����Ά�<�j��?>!�Mdˍɢ��f���بʏ�Sw��S��{l�Ri^�@�$�]��,�j�?*%���Tិ9}��D��A���5'����h,C<���i�>�z�L� ^f������%@oໂ�^Pw��'!TP�jl�����J�z����O�9��1�4��Ĉ�6`������� �O����S�V�j����ˮ�5�i������Q�ntm]GJ��$�Bھ1c���w��������� ^��W���6/o{&�����/���>�����2=v�#ޝF:�H+��@�fO��7�e�:�s�}����[�-�����%�N%��P��fE�z���J����Y0|!������XI���_<fe��յ����=Cz#(� ��q�'�ϒj�rݳ-�P����ٍ����ږ��z�<QQ�]?�ma����} �p���]$�"$��OOQZ���S�+��P�N�]���ST�������d�4��I�*���r�9���1�I�M�YM�9�$C���D�D���N ��!IXEB�S��jF6��o�qt(ό:���}?؏�#���?P�{2 >�8��j������Y:7�U�߮� 7�Lem��&��c	&C���oM�T�s*����������H�M���'��!�T_�0���7�Z���+��=R.&����20[�.�ߍ|��9��.؉-����}���*E��;��'��M�:��Q��i((�"#��K��~�MErNf1_ĳ��f����� �d8�+&�!��#\/)G��E<����gkt���B�7��,ov<*Ĩ ��y'&ʜD^��K(�%+�zgu!��E&Vk��$�G_{	�@Q��e�GXzO����� ۹��������$�Q���{
N횿�o��>Gl��*��ZF	:&��ݒrPW^]����;�p|�KWҴ#���ΘT��)��y?zqLi	�w�Bl��#GO��ѼYs%�}�������U�TJb<w�=i�s�^5q)�YM���ס>�wpz�܄ĕ믖�R5��f�7
	�~�J�s8�'��	���`�L��3^�����s�A�~eݰ���(ݖx�h�JLq��q������v~ '��s\��-Hι�T��=2����LZ��j���S��a���\���'�O��ǦZ�Oi�e��<١����Q(@O\�HF.b�TY/�rbno��]���x����T�ä��X��c4*��Yh��^M('P8��_C���k�����"g���L�/<�T��.�b�V���1���*�(]�S-�u뗦�<��O�l��1�`U$��!�,��i^�y�D�g34�k m-����e�󚯯5q�o��`�*,h�����;�����Q�&�vZ�4�([)���x�Dԋԝ^�5.�Pk�C~h)����,�+���4ӆ|^��O�0ճ�q�ū��'Wj�VM�+�~�maa�`��izfKE���Cyb<��5�i���2�#o"<|��%����zc,73�V��J߄�3���wq>��y{
bI���M)���7DZ&��B���I���+2���^To��O�>��b��~�g�A tC��U���r���:���O�B8R=G��iRH�?�aH)��EQ��&�T��,o�_q{g��M��7q�&r2Kb�,�Pʞ�1!4�Cn�I�d�6�!��;�d�-�&c��}�p��gB��g�Eg�i>?�c;�
\��V&�9,81�G,�R,���3s�hyN	�`�&��ܸ�>��9����v�b�R�zUV�ӧ}�̇�J�:5�+��j*G% b(���j��B��Y��T�#�$Hl�W �)R`^
4��UH���C���&L�%?Y:���B;�7q8p����u_F��n~��b�>ߣ[������.a�^T���W��d} q�;��c�k�1"��ʌ�O��pN� F���?�����&���w�VJ����ȨV�S��ڧD�R��bL?5FL�ިX�-,���45纮�5=���F��"h�	��j�Z��
~�׈y+?�~!m uq�3l���6ad?/�x*�����i�OBC�F<h9�1�Dsxd���"<ŏ��Zt:����)zp�a�	��5k��|@Х����Z`있�RX麙L���RC�^�B����d�E��U��CE�ۜ�H$B�i'۬X�Z�����"Ow#�s䅍�F{
����������_T�8�Ʋ�g]�Hs>6�&�a�jL��4M��t�j�
6BP��%	xT$��y��ǹ�%o���"�[��K��#�.�#�I\����sLs�׸�ٙbO�/ƇǗWU�?̫�s͔�=E&�J����vbJ�e�V��ԓ����.e�S�y��L�[
I���(o.�Qߝ�9B�.&�:p�@��n��p��b�
�8��[��ދ �)��齕���������������i��o.�`��iRr�n	Lt'��ǭ��|F+�����fC��-��]�P���s�7�
�:/�(��AL��1�u�Z��)NX��D	��p|S�g� �ca�O6��FP7_���
�N��LO�u�k��������q����c���w��hޭ��ؒ���n1J|Y+:��U��,R�)���V�b������)67��g��t$*��C��FZ�l:u�N�%�d��R���D���Y����<������*�i��V�mK��潣sKeh��l�%�Kq�Fۍ�н.<S��.��i�9t��ME��T�rVو4V��	a�����C?�*q��o�V�@!�!5�L=S�����>�b����4*tv��s���~J��
���u�Jh������	�d��ŋ�za�r�ԍdfZ��o��zp���Xw�4,�[r�J/�`����"�vt���c��)�O���������tp���i9�I}�z.؅jR�ȴ����fAn!���5:�7����Q��ˈ���ȕp��8=#��!�=q�U;�>/���N�/�#�k�+ü@��0��j�/���X>8��Z��*O���>�ߊ���~���dTt{u jt�+�tț�xܽX<cA!O�n>�e[�<{��u[�)9�g���Q����%�ٽ'�t��:�K�{�dPʮ�r�Cm^)g��:��'�r�_!$Xk�^�S+�0A�G��YA
�1g�����w�kk���1�ʑ㍛ӓ���$��Ŵ����tB�#�1�R�w����� ���W.��lŸ'!�����|�|9�% �>�̠���w��k�m^��VDr �ʼ�ua�%.��B��}"�%�Pf��z�(0���l���aq񲇃^�7b*�N�d}h	7�m��rP/��b�뽁�0ӟb�X�"��_@s;b���@���$��]#)c�r�1qT�)��*��Û�4r����ty}\��j=�x���d�bS�vT��W*GmS���[��pI\�~u���'����z��nx��R��B
��v�1[M�@T���*��~�x=�	c�yU)����_g7�~�	A��}i����ro͇R/w~d^u�>�KV� vw3"C.���{���I	�ˤW*܀
�9�n�'�MP�g���٩��/�}���qR>a���&��u��N�xV�di�A�R�,*�D�0_��m�q���n����uϖ<.��|�9>����;���U�N�\���":C�Ug�4�B��g�J9��H�Έ�*}wf�W��M��:�u�rW�?~/l���@Ό��P:'ЖT���������*j��Sx�S@�!�c;�3C�͹��E�
�Y���f���x�K���,�+\*aS�;A�f)�nD`Z��{Z>��g�{���2��E4j��EYƱ�-g�������]�r����p��,�L��.b�Uq��N(F��.'�T���St��as��5�O��l�w	H�S��e�ɨ�f�v��sdaٽ>�b�����Z��1���~�є����tLsa�����A,��N/nYa����BB�B"}�)��T2�{�d.����t�p�/��$��5��w�����n(�:oj��3�܍��])��ɳ��dL��XX	R�K:��uE�\�"?�)\HOS����=�-^��"�}ǩ�;���w%���ZQ+(�n�WQe�U�F�Mi�bX��F4���,D�q�E��͂=wR��Y�D���'q8x��i��-���n��aF#$�\� ��V/c��
����${񱹎WMf[k�r6�-��9ܕjw0O[�!���Q�����-k{��L*��H���C!��󆦱�7a{RP�a͍H|/��KGJ�j�fH)?+�������7��t�E4yq|`~Ծ�D��o����V��ؚG���2"ɷ���OVҚ�q��K^��B�a����^^�ϫ}����ƫ�n���U���R��iY9���N-$w��X�PC��M'����Zt����t܉+��g���9��N�x}����n<� ���uŝ)�,�@������b��~�ė�9��% �r�/�婳ځXa-|�\�l�g��%Ѓs�����u�g�c��0P�H�]�䗫��li���H�}5C�;���')1��AU?�۶9 �u�dǄ�̔�DIB �A3W<
v.�a���O�������V��B-��_�"�ڏ6��Uf�`�ey �V<,{��1��}���h5r�[�<=Xު�-x�v~r����c�$��cjQ\�X�Q��;��)/1�􅉷�^O��j℔���O,G�W�ʩ�f�Ý|F_�_<�<� 2�q�)�h��5z'����X��P<��F�>m�(�iU�����Q�^�xI<��PВ$�M�3�cT/�!�Z��겟�v����G�ܗFz��(ѱ^��S��-���[t�w�O�;[��t��r.��$�T�E�iyt�%��i�Kk$���f� �:���!�4���meg%i�N�F���Oӏy��hN��ZJo$�����D�+uԽ�~��3J��Q���Q�J�� Mw��"6JW����&>դ ��w�)nM~������A��%����`=��o���/���&�˴yb_�W��dAl�AVKiW�Djh�W�<\��� ���p`	�˺�/)�f��-��}����e���,q��ֶ��]�j�S7�G��$�Կh����/V �D������	����y���]���-�bq!�y)��-�u����#��l�ǈ>���T���#;�/p*�ͷ�T⢦j��"��9�ьE�0z��\�ު!��
=T�&M��ۦ5��e9e%Z]_L�k΁Z��o��y7�mQZj���;w���.Oe����<�;�G�q-��	�=w���$>K5�����M^�����pB0�2�5r�Sx=��Ʊ��,=N�?d��p�'�4Zɪ�J�r(�C���
d
�w#9W��3׳��o�4������ZN �&��� ����'�̪$&ڀ�	@�D�ďC�a��P9�4ʝ�Lt)FV�m��f�W��WdZ�kE<%>O3.םZ�L�� �E��Ϛf������l�crk�8���m!�PP����A�U�X�m�*�[�O,ҦMӥ���2l��y S�~U��U���j��ALD���"����潅~8 ����^�X��t@����+��-᰻�Xp�a>��HE��t��Ļ���P��A��,�콟u`w�-X"��(��{ZV���������cCq��S �:�^�4�>w�u}��(���Qΐ/�FZb��sq���ߴ��C�������LnKB�P	�(8��oYt�����4Y[@�����/:��xY��v��I%{ʉ�PYF���?�d��ބ��L��7�U�4�A����f��7�0ζRϿ4�	nE5:���4���Ã�0"��H��5��p���У�&�,�r!
��u*R�xB�w�)#/vq|I4��묾;{�ͤE|ʮ�ihe7Y�dN�/�
(KB��g���vj�ܝ�iP��+��ESb�(��N����ֲ�����\p!�X�m�����1�}���#��D� ����ʥ��f[1�rXJ5�"L�U{�(�����ź܄���S�ba����A��*l_.�AYho��A 6��Nl9������	��<uÃ���� �3�uS����R~�n/��;�F.g��%}���_Bu>��E�� n�
�%z�a8�vR���'��΍��<e��`J���O�Z��y(�{�HϿ���7�°.+.��Cr8-@L����eCBڵ��K��g�Z���Z�Z#�kA(�ێ'���Q����P�4��0E���9��RD�dp%#1��ҬK�%���R�����36X_M��U�`e�4�Rp�lLL�����!�||$U�îob���-� �$���~N��O�O�[R/�Hh�n (j�����3p�9��T��Q�X�g>�$�BB}6��C|a�"p�!�#		�|Ԡ<�q�0�����=��ݥ�~B��7����OV	��a�Fh���v��&����?���2����nÐ��K��)B��(�p�͸�m|;Yj$�su#�5MU�����C!�6\��!��0��9T ��s�O��zq^��h��ݽ�.�JLo���r��:��ç���Q{%�n�{hW,�JB���lB*.���8��Q\��Zx!�Ql�4|}"��da��cb0���Nhn��^%s�2��s��J�?	��P�tG�BE(6��$��ȁhE�$�(l�'�%���ӗ5�U���1�G	1�0Q���.�����S�rK���u���U�v��f�ǫCe=��?�IQ���s^A�����g�r�7�`U�n��	=Y&]�1v��
IݨB]�(�d���%���I�.6�7�K�@��_��3�2/��d�@�sH���%��w��,UAB��gL�sW��a0��r��R���/��]e��w��rɦ�!����"�D���l��Ad;oūft	ś��0��爕�YS:V�a������t8x^#�X�#���� �y��zfBEB�{����q������ ���J}���?�$�a�>�ǉ�Y?�Yk��o����r��$S�rk	���o۴�sz������q2y�D�H����~t��5��Ņ}���Z҃+�=��@H�=pH��[��-�?��T������8���_�`�FG�v9CGUK�����M~{䱏����x�����ܫ<*QW|��f󟲁漣Jr�̚���qU�f�a�<5i�=�]�Y��XCJF����f4����5}F�"� �,�{sTh�?,
�^@K���~2D�h�v������7��yE�&L6�vm׮TV�8�*)s$}/<E�F���n�fdvx&��3Ģ!1�V��8�8w�!Q�=�� ���"F?Q&���� Œа�Q��d��- O{�8��"�e�١$mI����؝�񚭦�2����f{��I9p︹���I6>S�,vI�.�jYG�7��-��2axվ��&}|��\i�J��w�Q�5�0o�q(�|f��^��/�lR13�ؿ/�ͨ	;$��p�7�������M�@��$Ʀޒ@v��O�ꉒ�J���9:_�Th�5�8Me	e-����%�\�2��v���Y���*7�	{�?��ߓ�$&���>*uA�Zd
|9ґ,��$-�U��(�l��-�K�S�=y���N�I� �q��֔�)'O�kɕ`X&�B��;��&�a���Z���>��a
���3�����#dSsdXrC;��L�����:	�����F�+:�z�/�Fze�*|�+M���j}L���G!��۰��ݴd�|�|���g���h4{�}��:��zۑ.n-{��[��eݹ�cu{S���UQ��t�^K�����S3��m��a��d�bCgSEPX=�ErI*���K��\dq�@\&:%G�7[ˬj�l���TE�E��G� Z�8�~I���#>�+��2���Ls��;���&ho��d�������*_�+�%FruC�Lgb�������fX�����W�+F�n��$��tRq�5r�J"���?���ZE�↮���NF/�NKvH����;��]�؂I��\�����MBi{����R��
��Iܞjo�\U�h�gPiiSC%��f��0;�qή�=,a� r��C���8��p���5�sM᥆��X�n0~07�V�@&3�hs�#~�-�N}��Zl��Eܦg%\�'�)�٦@%B/��r�M)�a]�p$Q��S����$C���#;xH=�{��F�ݱ�^@Q
V��[i�4���z����S�m; T�)���ޭ?�m�1,/n��;��Lt���>�d���`[�������QC��=��A���w&�\/�*6��qk�@�߂�Nf�?�B�z�!��t䯗q�)Y�}݅Y�&d
��>Ba�C'��A>���6�쀬�}_([�r�������h�q3	������v�k9�E�Y����*��kk��������Zڱ��e�g���)K�,3���y�K��*ϩ��$�7��J��9�����3Ebċ�����fXܸ*��%kE<���ۉ���cͽ���[#�[�H�z^���;��"���k�=��~�� ��%���r�6�٦�Qd�������i-�v��`^�,�5ZB(�X��`��woH!�����g����u��	-U��q���1���&��*]o��c�����DK�&��Y)��eG$��h.ی{�yq]~��{�`_�%�d��îrD�
=�ֶ��6��6��#|z	�x����T�oi}5�:c�]��ńPXk@�q�(5���	J]fA��F?�x���nE�'8A��IQz�p�C䔮%_P�y��uo���B!��)�W�v�,�z�	�m�ʖF�*.UAZ�`���Q4�JT�� J�~ˈ�M$Q^&�F��]��:��ܻ/7<(��6>�/��PVVZ��[~��@�zn��A%�N�P�ȸ:�r`�7b��0�ձ��i*|����腿�Beg��G�CI��.�-��hs�U+�:y��b�����1�R��-���c19���&��Q�$F5�jO�_�J��}?ax�!�_�r!����P/caPx�#ǀQk9{��)��#�y�� �Z��i?��n	��"��RA*�Vx҇�"�k~���'i�&�M��O�w�kޱJ���*� y�|7��)N{}[{��-�D��G�,û<a1��X�͊kwn<��h�\�����U.П��G�x6�����>C�w/Q��8�tf��َV2�伞�w�L9�7�JP!�-�M��_0�9��p�UU\+P+G��5��C�6 V+�\��%������d?;5��Y6�}K���)��T��m�E��w�����[��
�����oh���M[���<&���
�c���=����=�"�	m�涬�g�z׶
���}"-�U��`b9�j�s�|q�a�|�%�9�y��;22@ٮ�V�q���[�'��6S[�>�a�o��X^膱�9�DC�<U�7��,y��n��4+'4��	���8��<�&��NG����f��X��W	ݮ�,�y�1���xco$���&�Ɣ,��'�1�!?�aV0s_/ �x6���&j}uMg(�z�65��.�͹��\y�O��?s��IV��qk��8yOL�яy�_|��/p����E�S?����*����)�v���G�� �Y��.B=Y��\h�wr�B��'�/�i4DR�i~�V|e��u�}���Wv�)|5v���A.%ĕ�h���'/.�;N�r��!dʈ�I+�n�+ނ�? �ށ˥�0RL	\ӯ;;��R���/�9�3���a��]��߯=cej|�R��BѰ_���9������F�hD���,����P����A�f�h�.�[�W"�_��|BH��Ņ���<��@8__/bPg=���}�ɔ��R&��ex��_��+���O��L���
�02^́�L��]0X(^[��>.X{�2�:;���-��#�TU{RX(:��r���|�Oq-���?L�� ���
o���-�u��]�
�N��k�R�>��i���+���8S*���?���u\Fl��mh�T�(�S:̀��
�U�Ɔk�c��P��껡�^Sf�T$5Ψ=���D��z*K��N�q\9�"{5�$5`p����g;�!�MU1K�V��v�i 4�����LӡW>z�<=_c�P��8?7��ķ���h!t�
�K6�Όv��5��X�Sƍѵ� ��U��L�g�������=EQ���VE��(3$��L��I�� �����Zl/�-�?ʽ�2ו�fh�2�~������A$y�⳻�W�i��]���<}t��*ng��8 d��eYq�����Z\"�� u���s¹w�5��;)�.k���E��B����2/��K��'1�>�`e.㶋�lE�IeDQ���"�.<��L���-CMuV�4ɮ`UP{j��̳jWS_��S���|��Z�G5J�x�WFC��ٌ�e�<m 
�0}�]C�_MnO8>��g���12��
�C~�ٵ�v�N�m�o����3���[6�)A�nq�RZ�W�+J�/J�����m��M�F�H�����CuNq��~�дY8VQ/D�@�)s]�te�i*~pb��M�V��:��F�*���{�V�h>K�#�&Z�"�a�%�f�w��A�w���B껏��׳��I5;����l��[ۆ�lR���5
�;gH��b0�\�Y_ޜS`�eE�[�ie��H��c:s�6:�U��Y�`9�L�I�0��}��s�(
�o���~��
D��.�U�����X�4Р;��R�|&����� �� �����/~����P]����2/T��`r�>��0��#ؿ4C7N�T�.�h|�#�ś\�퀳� l`>?��Av��-H4:H�N]�^�y;%Ŭ⿋��Ch�1N���@�>������4@�I��Ы�"Ι)�,��{���_�ыGLmԖ9� ��xxR�m��/ۭN+��3�=T7�A�w�,=PL��� #Cf������:w���`�d�D�sz�����(�N�V=~�d��vzA���f����Z�-�/��pr���i����Ī-��LN.����u�U�
4�<Ep\����fӂz1��,��e�2�S/��ӑ�,�o_=�j�I�)��6�*ޫ�y�eM�QJlp��>��M�� !ՓN���'Pz��cf�v*	R�-�	z2��9�%[��ٰ��%�M'Y����cM_E��7j���N��`Qڥ�5Im����hR3P�	��k�e��1�d�eu�xN��x<i:TS ��%���{�Lb�&̫�3�L̰<�b��ѧ�r��Y�� o�__dr��_�eU_6nM6A��$�������2�c�3�EK���>���K��B��tH�?g�H߄��͎�nq��PL��_ޮ.�۴�QCr��|��y������8<9��d�8���<�����w����@�'�+�)A+�R�q���ך�˓K��W�B�WM*���IDQ�Q�S�.uDP<��`�}Q�M?�$اs���e}�%Y���~�%7AnP�$� �s`A0ژC�v�}S%�*�33�/��m4�A1�J_�����G���Ýr�d`� ��c���D��R�X�ʹ�]d*Mu[��g'j�=��-�䰯��8&I�Ѡ��d�6���J�6ȓj?	[�
w��*�-�ms���D��A���ʁ�<V!��x�{���E�f� v���ŧP�����Upò����h����xPGEV8��K�8�}��)���;��܃�-��/��%U�Yy���2���a6��9���XN��I��W:�9�X&��nY��\�{р, ������+ZՍ�{����0.�^�.�%�Z�Eh��&=�� ��N�8a��7^7�^����u7�T\�kl4]�C�sUYپJ��r ����|tf.��&i�2�����3m��i��ǥ�M˸�O�.t�bh(��L76S'j`F�u8>��g����%U.A8lLj���Uj-��L��r��i-!��� ���*a���s�#%�h�E�'�SiS�+���>��1;��m}�,Y��(�Oe��HU��+���B�g���IAO��s���k�֭����}^�S�%x��D�`�&�}�����Eٱ���!Ps��Z2�]�kq�g`�U�&�-h0�E�~QQ�Ų�ķ��s�_�k�������o_���X�lbG�)����50 5yyp	/$�|�e����6�����η�=�×��S_d��ֽ���1໱�T��F��!+�
�aɾ٩Ӗ�T�.�@E1-�p�ğ�zy娎��I��*c�%x��|e�3,o���	+j����I���.||2��7����P�f6b��x���Ǣ@h��%���!F�/ɜz�G��IhS�ɇ���h�����x*~�|�O���@�g�<v�&��{��7;��g;���9\�-t�:��.��l���x�S����o�o�F�'Nj�Y��Zo�)%�<&d�3�4A�u_�}3��=$^�%�cO���`?���.��n����M�~R/�q%�)4IKcV>��1�ׅ\zvI�0u�PQL�9H`��̽������LӺ�MU��Ƶ��D3�L
��fKMm��}�� �a��4����&�C�����>Y����*o�IL��5�:)E�=��t��df�[D>��0��s�~�(?�#�1pA~=X�9�	���0x�%)4���{���6s�ŵ���u�h���JAqMW�Ü�ŴU6����~H�VH�H���W9�
p��J% -Y�R��I����ϫ�'����O��L�R����ۜ�y�#~
�V���Q�%�pU���
_5H��gw ��k�C��c1���HM���� �j�$C澄�c@�� 
���leMH>
~�qj�^ J�Ѭ<&i��ݎ�џ��?�~��o�]�g��oC���VU �J�f�Y�����a���N��q�_N�E�����9�p.��І-��X���on�s�K��3�Q�����R�`Ы�	�k䙮���E*��CUQ#��J��F�%W$p���TQҗճ��!l���靊��]'���t�~RQ�D��ę����o��\�FH����6��P�K�#ؙ��,9��rb���]tBz�l?�����C�W���:��6�/#!ZF㮜y��
O��pA�t����pxJȺ�=$��(������G��N�+�$�\�>�N��;�z[�A���J���>v���6ݓ�Q����C��t��C��X�6�>�x��s�F�Z_���^��7�RM�L�H�F.-F�(Z�=K��;!�W�!/�^�EPd�Ur�Q�(,�{�<�a[��%�%��3D�B�̉�������C�ʌ�Us^����F Uu�wi�'9��уe�b�]�J��ki���]�~�V$�y�����"�(��J��_EDPZ@`=�u�H:n�T�c��߾}����[��Oj�\�+�ID�	�#�`C;�3_�f�m�嗝�0,1<G�<�r�}L��ZLaN|�a�B�F�.�V��78��!l���+���u�H��n�C`�`� #@�L~����XG��&�&U��FȚj`>�/i@T@MV�/'K�N�8d�yE�ս�BbZJ�fr6`oڕZe�R�9A�=���3�����/b���^��.�ײ��n#X ��8rj��A_�H5�u�`'�.L���u�RL�����kM��\� WT�ӿ�̷��E����I���)��da��:��M�h�*s���j�]b-������%B�7�c����{a@/ύL�-x�-��W�b��wN�]��H�۬2�4���:���C��< �T�����ؼo�~��@�+�4��>Vp����>k�eS aa�I��p*�unc3�����1�V Ua�K�3�+�p�bz�h�Vmq:��ksP���H�	]x����m��~�p�Dt�{<W�k��*���_��=����8Q�{ɕ[rnhn�n�y,�C��1߳��ցc�3	.[��"Z���yU`��*ۏ�p��'L�N��v�;���y�4���_ �]cl6���N_�	:t��(\�	�� �@嶱U�q��-������27� 1漎ܽ�����y�MN��e�"���E��f��)@��0 ��)��Y��[�أt���I{�_�Z��df�(���^�'�Ø5��o�a�	�]�m�}�������e���^H��*�W�"�G#�S�~��������.0�����19�N��� ^�"�3E�K�kO�_�f=�TR/�P}�mO��0&����%�4#�2�x��6:�6��PU�t��B�k�����ܖ����L�	�/�0J��ô`@<��_��5@_�:Cfv9$-�J�Em!��Z�6b�\u���@@¯���;��-������]v	ۚÁ=���{�t0;�j T���tπ��8��������1���ܾ�7r�m��_"#g�Y�::ix�`B1�]dyL�P��"��~PZ#�'��
}�R��Ù0��!�Hһ�<�SD-�bX�_�5߇�s���^�����Z���漇�$���(*�h̸f�����@a��Y6�Y$�N�a��`��ӃƐ��^.ѭk?��(_Ч����({LK18�
���X�-�M��i�C:�͝M�uVxN��a*�-54�)qne�_�*t\u��'�n_2j�~��]Y�.���X���	,K��\ѶwB���_��G%q� L���6�x�k���Sv���$��49�gV~u������XB��C�{��΅ae٤^u=#��/f[�C�����" =j����h��b�����L+����!Q��M�$FCi��/Ҵ�1�!�V8��yh�_|�z��@=�.�>��4��V���w
�6�	C�(��ʭ��N�׈���&3�~ǪW^=�Tꮡ/"X��^O"��҃�Y@-��ih��1���@�R�2��`[�y�>Ӱh�Z��8a�Hi|0۶s����Ce0GF�Q����L�����"q��'�ܑ�a��t��QNR/�4��gD��ʷ��f����ە  �T-�89̈́BS���%����"��K���(�RáMу�jx�1�\�c���p�oS�7?(��b�$}��r�I͗�\��"3l �xV�8����S���oƢ��Ҍ�}Ue�NW�!�ۈ�!H�8|>,5�.)����L Fӭ�/R�J��#�y�?v«F�q��R�G>KJ�l�p��oV�g���ݛkC���C#��F�<~lJ�]3���,�h�t��������I�ʫ_ ߩm�SҤ�n7�G�*�j}��0)�<�#�5#>#%q烚��;�v��"',W0�`xF,��p��ӂ�`}�XwM�uT(��L��*9�c$��F{G�$n�N�y����j<���&�#����{�FG����S��R @�r��}51�)2p�#�(������`�zH�p�ؖj!j������jB�͞�u�)W\Li�Rw�#�s؀rr,Ap.��"%G��������(i���x	�����R��R:d:�WG�	�ߏY�
��F7(I'�U��x�w���C$������tW�as�k�k>�8�zgi�U� �& gN���'w7,am�H��Z`������	~�L�ԍ4�_c����D��  (MBu�q6T�P��yr7�-K�^�y��{����!l}�(!�U�s��tG���!�%�n�#�tW
�����ܲ�`��ЊB0�GW�~|]��$NG�u���$�&<��͊:�7.]֔�u��}Y�w����O�]�o����*~X�jux�'���z�Oo%p?���1��k�O�@��
[_�Z�O����U+୵�D�@_��s�Pv�k�ne1���D�hq��j��;���{o�<=��/����|H<�|�ظ� �z�6tq�>~��e�M��u�Q��PigY\3!�+�lx��	�Mg���-��U�ڊI��5W��XbyIR� y@�`��9'�%/��8���)�%:6���%Ɍ�
�p7cq4S�Mܰ�p�_!0�K��}&�j�7(/���#�b����~D��9��*�9g��D��id�l�U���<��6[�)ZK�H+��[�Q�ے(����#���� ���`Xpck�dv��l��{�U�jM���Ms����{s�t�� � �1��)��|�H�m��N���]�"��N�!G�3��W�_�_.�w �8]��*[8���b��^k���V\���C�w(/S 	��)����� :3�9�J%�~7:[@hH��p�?HG`��k����� �*7`/A�u�A��^��a2L|��̝�si�#v-�~��z��4�eg��ww$A�ۀ�M ��^\UwS�K�q^��:� 5��$����S���v�����7�?*�%�z�r�m�6	]�#��v�!g>o���a�B�RjL��t�&F-�����`�ΊbY'�w<��t��^��;��R@�m�Æ�d:�ߞ�_?�u�ٜM��R�Yɺُ�NV�O�_�:�$J��汤�*�Q!#�]��KE��8�H�B.����c���L�!��/�".յi���s[�"EK3���љ-Uu}���	��á��4���5��u���|kQulD*2]����Q���lcФ�[ǀ�Oj0���zB�R����kS0�M�h-@�"^��.mq��	X��9�/|��Gk�ep���[�M�x�Gg!�@��������x���| Dli�a ^��O�p^�4�����NGP�a��D��͏����'��9G��!!,+#���U���(��hwګ���I��s�x�TWWE��"����x�lc�,�Z�����]F��W�"�/����'`f.qw�5�W��*�#�pd	�P�U��ZA8$��_q26$�:�4�7q3�ȭ�Y㡷�~��u���EG�0h��$o����q��S[XU?�RD��\ڻ#V�v/)t�G��)�/��Aq����I ��4��MUBha4�*��W~WQ�����n>A{�J����`K�m)m�<"��c�w̢�t�I�s�tB�0J���ɜf߷c̫�[�V���<������q9/��Ņ:�3��J���okq��+u\^aI�?QL��3�A<�Q���U�y��{Ncu3‡5JKzv7뾱5�.�3U[\��9�`�a�
�Fs>:��.%��Yx�IQB��+�%P�f�[�tc��n��q�
��f������-���e�J�]s�)C��xRQZ�M��{(6�h>��c.T��P���C�[�+=�9��mCS�i����T
֡���I��a�<J�\<H����J���� �G&���,�-ࣻ�9�0���"�����ܶ��s{�S�x� #I���Q8i�����g���":3��?Z�yb��CUS� F�,�=�Yf௽��k�ǕgX�g�o��˫f�?�ȟ�Kp�%�� ��@��<Z��������k�%l�]��R�˒��<�?�I���k46�(��,�*@�)i0�0D_�*xzj�9�F�!�'M����}f��ڦ=rvX/�+,�Xv�(�eM�:IpAS��`� �m�>�I�I7��'�G�ڨhZI��h�Ґs�;@V�BA�a �,S��L$�H%)H#��M���?N��/m��0��Ǳs���6��,տ��U9T���'�~Hv����:4	��%���D�qP|���]¶�l��%4��[�0cݑ\Ʋ,�)�ib����,G���_��.�g�u�sw�AC/CZ2i�/	��;6�7�z�@[�bK�)����Ⱥ	{`h�	w�M螈�ӆ9��� Ȕz������ʼ�QE1��F�2�GSMA��Þ�Tw/�A��uǧ�����rR���u`�ݦ�u�꾻��\c��Ƽ�`���	g�����K���.�sS�z�^J@����m5g�����FwÊ�%�&��Fg��B=?�!��x�Zy��e���mM�B>bi=TҥA�X�j�<�Kh�9ʹ���9Q�Q����u�se��6�L����՗�T�\�Vgҕ�.Z����YI����zQ�Y@�����޿89�6q7�f��������R��sF�����_;�u�W��&E��P�^��z;�߬��Z_��>�jю��`юG�Iʀk>EK�ƏI1�3��8JE����kٸM��H{�?G��~�	����aF�p�0��@X�1d�����M�{l珔2�� I��pL�x�[���Ψ����w?�xn�}[��7�8Ѭ���GL�@g}��,��xsu�M��\�,�h�K%*r�&���y����iř�o)WTB�v��{rŝ�� \,����.����&�b�;��%�xX�\��)U���Aud�L�q<i}�s_6�9JB۳�/���h�\1�r0Pf�Z��y��j�@����FN�/Aӎ�إR�3�ni�?�_ԉ�.*2��w�]����~i�q��gW�+1�-�'��0��
z"�$�0&0�v�.��L���7d�N�Mfe<��!�BƗ�{Z��C t��m}����+i��#.�E.�G���Mͥ�����FE
�S���½�̩�����ɍ�.����m��UK�Q�Uһ����3�7��Y�Mw���4�f�f7���;3�`�_zT�Z�QY-%2C����D�TQ��B��kc�驃]�����OWZ�n��m��	�e�"ӡ���_���'P3Z�١����ʚ��V�un&�� P��<;_�K���`W��2H+FLjP
�i�v�)�j�q��/vHN�!�y�Ư�sY�p�X#��O�#CM]C�&�RCvC�	�T-x�/i�z)������v�lZ��V�d��
�.�&�'	�A�����^�E�v��Ŝ��O߿�i���0ג*g�![1ڄs9�w���f�9��7Xcxc����-�V�� 4\�B�[!7��N���K�!���s����� �쁥[�rΤ�d�\�a�^�+���Ƿ�f8����A�kb72��hh�x�9�\�%sYo�f{@���B_��M�D;�rǢ|TФobw	P��AM��cBa�u���8('�&��;Ch���<�(Uae��|Ȭy�{���O�2ʯ��DAH���y�*�e��ѓ���0�\K�}W1���#�0�;reVI�5�E�5*�[^�s@��q�SR�+��-��r��^q���ؖ�� �L�ΰ��Oy�!���.���>�s�DzȪV6vC����ety(���C�s�Ո-n��՟�)���§c���q�!�@Ѯ�xU��Ķ
,6�Ƣ�n�)l*��W'Fo0�!S�i7��L���O����/��}(����PM�$B�[��T̀iG��4]\<�+Qj����`<�q��N�L��Eo��7U��S��0%mɝ���h�c�O폜G��3:8	�'��y0�r��h�X�����j�5eA�
y�0�_�:���#�.�Y�rh�rq��͕�&��� d��br��=Gf�૮�����/ȶb@��J�%���OzP~����9&r�&G�*����A�U�ROzS2�y�ų�~ǻUoiA��)�qS�w��G���g�(�ZUkx���ᒛ�d��z2�8�m "(≃�@Nw٪�N��iI/��
G%Mkn����z����(c�B:���y��#��u����Gsdճ��}�!��wX����k������B*$A7-�,B��P Z�`��Vx�D>f��sx%Tr���w)kf���x 3^Hc2���r|6�AzD��s�ŏ�ښB�>*1�З��q$���(А=ӗ	\�&�3+XZ���VE�
��(%L9�̯��z;!ԛ�-{���`��g2���n����v�/ܙ\��g5)�FкY$��h�ek)`�C��V���r�$�+.4=}�V������.�n�f
%��W��Z��o��(z��b���\�qU׆D�.���5��#u�4��k�Z{�k%��`Fo��<ڹΡ�N6��a���j��v�P��=g�ßL.��K��Ɛ��|�}�CpAXj�~p���U��3c.��"�&�y����X'����
7�A�d�I�m��uSC?�p50QT�s���)�n��c�|��TO�4�6:�'|��E��
�f��vr�&yL����0e�)+�0�qג�mu?G���v�7�E$���K�j�]����F5�	w	�*`�"a;�.�������a��H5Z�`�`j�>J�s�Ҳ�x "��g�CK�S +)��l��L�:���V���Bްx�Ҿ��>K=� ������� T��T�;r���=�"2�U�l���a�x�s���h��t�y�1��O ��s��e���|�J'���;~L}u4�L�4�/ 9ZN>ѷ�c���D�V��*rJD���_��Z��`>=�M�
ѓ}���G�Ɖ�x9�X�>�ښ(&l�=�P{�<�^�ү��j�a���P��6��NQ��yh��e�r�6|�����:Z�Eo2&R�P�g)��J����)Uw��mA�q�%$��D^�&eΖ��r�ўϐf��]�7��3�t���KY6ߏJ�^>�atdK�r�����[w�`���\F�dy�}����I�v��f	� �@���+�SG�]��Z�=�ο�s���4ʬ-�wX���O+e��!�{��R5S�:�����e�NMc�(]�2�&�@�`�(v,��+�d�(��Ǩ���o)��o-u��Y����A�W7n�� �u��u�Myh(�ī�F����'},,޿�۩i�Q�(54�ML��T|n��fv.�-�7��e�t�P�d��_�ﴮԠ�+P�2��[!F��@o���ΆR(өQ�W����
�����0�L��!����lg�����j�u�#��꘻_�b���̸x�*�o�Rp_4?�v�����r�(�+,�2~3�F���7nWh�zA	-?�O��n!+(RԷ
&'�GQ�V.2�oܗ���)<����c���4E[�{=��)���!���_,���@l�+ξ�q��}�WRd�� c[��gK�=�>E��3�?�����3:�<���g`q
eȅ�D�-8��o���5�÷��3E@X'*��G\
����H4F���;<�7�J��يHxyZ�Ys�P�A1��&0��E%�|��u?�[b�&�����H!��
��%8�{w�.�,
_��C�7�ۏ?�����@3���P檦W�����,�0���k<X�\�GsH�ܽ���[6;���1M6���7�es��V90Cx�D��ePB��'*O�a샊*w4��N����äW}c��b���#�<���\x�U-~���$�c)��t��s�%w���f�a�g��jV�i#�.����L�[�=�ob���-��D+�1�d�>R��7n3����A8�bo���n���v�� x�٤�h�z59��\x'$'��P�X�k�Gw�$e�R�y�,��x� ��u�B)���X!^�صd
l��N�η�lsL��5ͺ��-=ı.x��ع��˟�D+SŴI�ߜơ�� �!e�W�F|00�(*2Մ��T����y3#�͠���#3BB��A;�����1��T,%(
�0#1����!~m۹R9��ˇ��)�υMG�W�c�_�*�o~�Q�kJ�W�l �y~��='-f�~�������(w_Y+��z6�Ā���#�"h�2�qȸ���;�!�
ֆOl�_��zw`]�HG�Q�;�e��$A��j��P�K� ���9RK$Q@�N�jr��	T��h61|�U7A!�Ǡj�%oc�eB�%7$��.���~̀�P�	�$�%��[.Ue�tþl|����o#а-Y�ckB�gt�+&�`��)U*u�?�n��~: ��,�L�<�`� J�� T �%0-�>;+�I@�f��| �=���zQ�� �M�`���>�����)�Ж Nߐ�%�sɕ2��/����U��ڟ(���%?`���r��9B
	κ�~�PtS��g���^ŵ���Aᔘ����O�,����*���9�e�5�p�4�P�t�?�K}�#n8)�W1y���
,��`���'��Ҧ�吚]z2�x08�:�����>s�=�"m	Î�锈��j��H�����~t6Ty_����:�N�o��������4@�+?4 !c�ΘE����l�r {����_����=	���w���H3��o��b�-��C��`���w��<S#�kj�����!|w"�� V�����C6z{��A| ���=/�}�%�F�·���+�&�d����Ֆ���9�(�MKx3��3��@�4@U|ׂK>�F�;Hl=�7���n����e(�7�@�T��'��{g
jJe�%0�)����H�b��\�H�\�y�gn�͎�7�^��"t��\���{c�&�U.ɠ$[�׵Ԉ���	�wlFP��P��S�X ��:w ������.v�`+o�ȡ�m���w���,����S�wD�p�6�p&��	{���h/�AԿ?~^ ��D�O�K>|$��9'(i��ٳ:�Hz�3���g\���MvF�ʡ��t��4����\I�>F C�)l���J���jÑ8�qO������֡"�1n��Fl�~��t[����S���͠M��N��R�W��Mx�o�F]�K�����r��9{	�dG�c��B���]�����a5��bRۨNTC�_���xR"��K��	l��ې(P%ϙ/=8��׃��w����+�0!NQ��U8C �k���o�)s�ه���Ջ^sy"��b���=�^��*iԻ�c&�d��y8.<2����Uƹ�@�:�9QP��k�1bj���%�ZH;T��~y�ߋzFh�œ���#ٷM���x8�_�Uf�7�Dۤ8Dr����9��J�?�(�6�\>�9����C2K�k�����]��ˍ�<�=���ާ��ȯ�U�XܑcP�7�X�5E5{�$��Y�>����
�JMRi���7�r-��\���Z���or��5�0g�̆�`�d9^ּ�?��Y������d!��2T�	Zwf`6W�n��'��0�.i�48yD�;����S���je:�d3�0`4r�T�*dh��^╺*em�l������B�ͻ�R>�D�ÆS�̎
�+�?(D�������1xw�~�������)�������1��w�3,�<]�:�20 �}6��w�勛��79�&��:����_C��[O��d�k�_0�l�����d��q�~����^������Ot��9��O�i�y���?@*0hQ��֕X���B8��@90Qv(��Ih
�+��P�_/��X�L @#�F�K<CsH���!�16b�lg]��a`1m��k�ЃBŎ�:��qv��|u��Ӗ�Y��Į�Ef�:��6����`�����L+�g���Dd+��H��.MH�3+]؊����Ej��:eZC9��
�w�!��u�t_Q�5ڛ���O��mbw��cEU�#��yܬ�Zd�J���H]w�[���M�)A!�e�Zt�Ê��F O�J"�9�:�r���z4Zu�Ƀ$�ƿ�^�o�Y��d��z�Ɯ0h�6�A;�ˌ�$�5ZG�}��ЮW����Y�Z���v���� u3����{S���7�#H��S�3�U�c���`�d��4�/�s��0�=W%EXGL���ί�P ��X�7
��5����/g��K���n��|̫,���Q���a�[b����s)
S��h�?t$�����(�������]�D�4�a�^�_��>˥���+ר�f?�zْj6U䱱 ̴�'Ӆp�d��d+��B�_H,��:c[l}i�P�r�t�U=K=E�U,�U5-6��9�$9�[ā_�Df"N�K��jǎB�*��6�`K�*l;������k�2��f�A�W�� �=A�{���fHE�J�E�`�pi�U��3�����CFl[��/��P�E]eq[��6�s�ee?=!���O�a���_�M�q��(�p!eh�փ漇<.��{m���\��'�`��`�_ɑ|3/7��Wh�V�z�I�Qr�

ML�;cڠ��1&>5C`M�\	"��mը�_A��	�o���]IQŧ4v+ k��"�{�=	�����8_���Z�pL�%���	�w 3<<���}���|�����ҳ�^�$vd����n�|�F�_�xi֢,W���KW��$��r��%����ZY�Ȥ�X�\�^��i�6�;s�-�����6 ]$���B]dxV�!�븤g��h�o6M�7'�Y��{wL񭄺rȖe��ϒ���� �w�B�:Ὺ�U��yA���5�W�|��g��t����#���9�ٷS�U�j�1j��V�*��<N����/�itz Ӹ�:����1����T���i�7�G%��Ol�4����H�`�W��!X}��V$�����.��VH��Ȩ�4F�ׇ��+�z��3
�{x��)x;���R��z.
{����:�3���P���){��ǽ	+5�1*0;DX���:9ԒZ� z�=�av�G�L)�g��|�qg[<Xa�?���o���a3�(��~�d꽴H�`SZ%��֭.`J�e���޽�3�#!�(ﻎ{�H2��ǅ�Rw|��ϵ���/���r�b�
��V��d����6DZii<H�_~u;���*�9��tpW��ϸ�֯�c�Ȏ��SF���<���$Rr�����u�瞖\c:47.4~��ht���Լ��*�-Z����e<7��:"[��T��ㄳ�!
"�1G3�Ù�hv!L˅��}-��<T�1Hu�5��$ ��NS�M�Rp�0�C���7��˧��Mnw�����A^��d�7W�_u3�ҍ�OR�)]ވ�s�IRN��Q>|�=s"p!�U�5
���b��؁G�.Į�Pu���|��ѱ�ߩ`��)7��}��$'ט.�C����igM#��E?%��a��!�a�����i���$�RAٝ>��)%#ؼ	|��Y�~���	�3)(�3(J��N`7���J�g�%��`u���m4��$���.4TEEZ�KQwS6��V�Bk�1zb���$�2�����k����:�@[�z���zTbU��BNi�&�5(��:A��+���e����2���<g`?��s"b��C�妸��O�4]�S��U�fL��ڶO��`���7v�ͨ�Uk�o���;�uV-�(_v���L�� >��▥d=�>�rԘ�_��$`�G�����'�>D�HH�,�~�nߞH	:���G0�qT2����A��+=�`��Z껌/��}g�b;��EY-���k;��rs�r���P�.�T,y0���"�O��^/��5�s?��#e6]�����!
�(�U�I7Dt���.��a�7�z�e�ȕ���î�u�0�}i�H[�v���wY��9Y$%/9�"TR+ �|8�N��S����8&�A9�9�mY ���.���������x�P�n�y��D�
c�z��|�d������.N>q'P�����2W�z������Lʄ	_��ݼ�{b����n���	%ǩl�9<Ůq�̌��+�
��nC0����(��	1@4?��d
B!|��s�;����[�p|��\CWKp�{/NH��?�B��K#RJ\�C:��-R|-P&
JD�!��$��-�%y,���8�V��=B,��^ul��y�l��̧HM7��_�͟��N���u�1s�D��a�tn_)(��`�P;!r�7�.�X�l���R<B8�������$�2�o,˵�q���.!��/�#T8~L��;�����)n���a�i3R
S?Eߙr��v�uj�_�%b ��)T�b���+끂j^-u��5����hs$��� �}!?��+4jO�?�K�tΚG����T���>[������q	�Fd�I�"�r�l���Ըx�.I���h�]w�j����V�>�9J�*�A�O�����#Չt�-6�=R*%R�{@�౉��EUQG�
={�Me��l�Z�:^�(C�_.��Y�q28xm5��MMjY���g�R�]@8����;��4�Ѕ�UR��� ��v�3��5R�Ǽ��P������~L�0�t#�z��0p3��ň�۞~U�ٺ����QC��7"���G�j)֪0`МI�rc$�e���h����5N��2�7ɬ&����!���Ly�	fBc�D)6�g��[�*��R��)*�b>��Mt���"���'�����E��0	�+_�,D����b����9�ؗ��r�3n�A�G�O^K��Kn�\b>7O}�L��4#էIz�8�%��61�<}I�3I�+�Rep��� 8A����?�6���K����M���4��_����,sV�|7��V'[:̵ڑ�Gh��L(�,ȵ����ɭ�}"�{��r���k�8�y8<�<V�����-z��Pr
&b��.���CE/!�6n'A��÷�&�%S3�lN���)9!��K�^r�}}
"��5�P�j�2��9b*ٰ-"0��sN�րDP���С��LV�k�˧}�zv8_��"�m�ǵ����D*	�D�Ah��R�m�%+2UA�ԫ-��9�"bv���\)�W4��x#
�Z����_�YuKy
s�g"�o��D,߷�W噍ef[�ɞK�)ɪ.�w�x�b��\(�����֜�T˙Ҷhiog�c�x�������1ƅuݜ��w�)�=�D��U��������l1swH^���'ق]a�bv-E����Ӣu�6>�bWb���xs/�qd!�Z�#�x0�� �N���|���*|���E�!�([u��[�ȹ��Ymu��=S:al�HDBb�i	��֜�e��\�LT.4�9�
���30^��'��v<\�� ���]�sqI��D]�8kV�"��/<�0@�	�I��f��&�U��%��$/P�Gh�5��]��i	9�;ɰڙ�a	g��9���Z�|��d��g�$�.��}�*'�!W�O61~f�`��ж�Ro����u� �5~�aڭ��E�qt���io��<�w�d�ޣ����{�x�#�S�!K7��1iU��⎅=��[y�(|�x�Tw_K��}UA����h�� B��#�c��o�ۧ�A�w��8{c���	�Ś�{>=���s��/gd ��xD���=Z�h/JQ�u����/&�kub;t���VbRo(��빣���5���L�
�#\�|E�(�3��"�q��Gq�T��̳�K.)���&�N����:]������մJv�T����\��@�hk�1��.�$�S���9o�Ω�,�U�2���a�]~>o�>��_O���g�����"�����X��
��N��p ���D0$���}�����z�<�ٝћ����^�/(n�3��N�L2m�|�t3 ���ɭ�*D`�2<�ۃ�`�TMܽ�:��u�4Kg�WT�#$� ��][n �4@�it�t�^�7�6��Lpa'��e;l%޳1�
ټ��{���ԧp+Ь�����s1~������rqm�k@A��R����Aљ~^���fzxa���� ��u6�(%�e��(��I�����F�M��~���Is�-f{��$]dL�b����u���1~S�ͱt7�y��AN���*���o�;��J��+�tx!��-f�u2��	��0Z]�噤�\s��ȵ@���l㐭������gg�5���o̜zZ����Xl�`��0w�?s���f�1_��,Uc`�'i�D�$��:9C�G��:T4�]?�#1�Ϛ�=`�;�e��ص]����֑9c^91��<\L�Ϝ��Y�C�%��šk=$�L�D,<�C�Z�t8��}�{��@s^���&���B�� AnbT.�E�X��đwfX�c�����?g+��g��"��Ϲ���P�~9��B+RnO#��0�e��|��Dٯ�L����E坮���}�<ϠNJ}t���y>˾�;}�&��5 �p�f�eUm���Ol|[nNt�
�q�1H=vT��*�
;��&��dN�pc�藍��{�5���6�
����(5
`��w�	�����|�bl T�]�C�2�WB�tU>rF����wH�� '3�Í۳���n#�� �)ӆ�R���c���eq֠�*��8�M������s�D)yʗ�߁h	�������1�q���iIL4oz7v� ���b���6�H�h��؁(�Pg���銱��hrي���@nE���&7�F��G� Mtm���q�k�� u�F��+�djdxLÓ�1ݪ��g��I3 ��U�{�g�������93�76	Й��%���&����Q*;W�1r�kp��]�=IOȃh�,]D�cMM��.B~�*/�Sk^�w�`5���¢��/��Wz���0-� �RY|S� &kQ�06�*aa2X�4Պ�/���&�1�\��|��!-�[eA�j�z��x��_�S����H~|�$ڽř�kϩ�S�C}91��iFx�t�
!1�4e���]�O�?`+>rZ9�dfm���_���qy8!�;+�T���sP��/q���,�wF6D��W|�I/��ApR��� ���-ޝ�S�!V�Ш,�!.���M4������@[��،�S���
:!���j�v�)���:�Q炝����{|�_/�ਸ਼��]9�����r�����@�	�Ѡ��ƈ\��`)n�������t�����CA�O�d���Ǹ|����z�	�\���
mFf�,�a�zK"s�2ץ��fKLě+*��8@s�]�h;��U��)�K{+�ޥ��?q7̷�Y��.આ��8��R��aa��h\,���!�z��l.�t}l�������G1~�?��yH��:�%��'Ij'���$�kM�5���ѱC�5���jθ��	��}�vx�1a�wq[rx���d��.1����Tȳ������^
��7�1.tb�t¾�G�`�Z���	2��U��F��f����婁$
�F?��2ݮ����,yĔx`��۹�YK��:4����������t���o����?��m# ��a"�iZ�� ���w��A�<7\����\���_������TVf���$��
��G_����xz����f%;)Jubàa�J�6E��7c}������hP�fL(/
�#�,p&�_��W����IA �Ͳ���?���lİ9��}<�w��ʇ���MԀa�䛯I�lj�k�*�nȳ\��>�=tx��Ά����u����M�P��7>�؋^���ث���-���� >(ξ;2� ��'�)��(�W7�X�[��8����Thg�'α��2`%3���*���i�ӘS��i�'[��[q|�JL��>8�����׻��h��S�ҰP��\}��r��L+8$�h�o�SS��b���	���1�&�[��mU����� �d�����A	Hd���jy�i3ǤQ������8.�2�v�Tե�Jh���>�G`؀��}���Y�\�+�:)���,`0����l�����?��G
+����~ʑ1��Hg�4�;7��n���(���fa�s�%76�~�YA}�NQG���*}�bY�'ê����X��YS(%d�K1��|8��Y�C�a��d��Xt>�E���r*���Dh�c�wZ�0t��˷oW�Y���aV����|щ+;�-YU'�t7�
�L񙡊z;�QRhJ�Xe����J	t�|��j���g�U���L�	��)�gR��X��[t��򅦌Ŋ�R������o�E �>ܡ����u@�H+�	�U�%!ɯ^�讅����X���Q�w(��, 3�RS�M�������w��ǉ�,rbR��G��ky�24��zY7�����C��D���ژо�@�n�N�"�檽�!�z̯��%�N��:3^�۵��
3���d�I_ݱ��E���r�A#5��(}[kڙ�h����2�5;̙4��	�.�Ԗ�v���"�L��p�׳W�Je�s+r(k�18Y���U�Sؿ*����P��bNM��͖q��4�$@�]2
���P[=�����0w�h���M�B1�e ��j��sh�k�K����W�W��� �6�%��Q�<�Ɣ�cD3*,�kn�'�嬯���=�hz��Qp�
���駮�;it�Y"Սl�	3�w��@�.��'����:hx@�@�ߤw8��*�
�{����P�ۑ���ax�҂ P�=4�.��=9¿��q;�NJݐ��6�b̠�A;�<��4=w��̮�p�uh�����ܞ}.��Į6�����b�B�d�� ��)����������}:�FC�m�kC���u�j:p��>�"*�J�o(�'�3s�Uv,���I.Z���sD6s}�}�{hƽ�"̓�ab��fW	�;
[�v��]�cx��P�ܗQ#���ya�2�|�`�	!m2�:� a��/y�Aw�"]i ���gh�����*F�|���I�wq��J�B�[�?��m��n�Wo���C�azTSp�Hb0�U-��f_q��8��o$9߁�g�����!J�1�@��v��k�F���G�8jw%��\X�N]C�ΐW�H%�O1_�lf~��B�c�O�O^[Y�v�cà�A�A{�Fo^*N �%[s��b��H�I��<���5৶$6&G���a��	�a]��v�9"�^�w
ҩ*�XX�����:���[������z���:0�ɇ2/�H�j�� ���"b��vJQ�;��:�P�ˀ�Xb9ƽb��n��=��<�����E��-��D5�p�E��9v^�:�'yL���U'S�0��[-��k�fE/��0��YZ���?�� �w�6���1p��������]���e��XE}�j�.�؟~���F��$����I?����G�_I(O�:�"���[[����vX����?���-��0�#)P��BS��@�8�,�\�������Ey��S�x�W�+;l�+�a��;8�����\..x;M� �O���_m�����,!��N&��4q���s����\�ظi��xg��CL��*]Yf�g��;S2�d���;F���-�c��׉Y�_E2��;~��k7ct��R��j)L'��-P�cm�4�5�FBź��	
 ���t��ֵK�#��ꑳKV\޵o�q�T��qq� _�n����<X�����Űo���;�)�QO:�+��?\x��u�e�۾C쨦E
�mXq2,��֘����(Fg[5��֘�l����5�J�z�,jx)#!���w��4h=�,��Q�
95�B�B�[S�vB����ۍ{����'/�uM���}h CA���{f����mT]���^&�S� �(8#5�z8r��\R������a�$�s�s��$Ȗ��GT�A5�6D�~<��ꊴ��!gPn8�7�Ki��}�7{lU_��ؐ����S�!B�� ow�jYs0���H3��B��`�s�C� ��|�w'�}{��������x��߃��!�R�]$�"�ց�UЉ�{�sf,ř�3��zw�H�O�t���vƃ>�#�����_��Zk��iH#Hfn���V,b������}�Z�c��"g�~zIY�f�P��p��&Y*��29?`������h6F�0S1|��M.i�W�eB���;��3q7f�O�dҟ��>qI_K��@��������t�P���P���޿tO<S~�Rn����en��!Ӭx�o�U�K����Ɍ)�j���
v�W6�yA�Q�=}�ujY�[��S��L�.���b����D��Z�����S�ܒW.��r}�-�z'��T'�h��o�kQ�k� � �Fh��Y����|��jΆ�-Ω��)����2;\�5�_�[�&C�xC�t�н�>�6�,29ͳ��$�5���K&�~m[�OdWu�`�+"�;N|�ȥ��:�ώ�ONpj�{��d�*;-J9�
?$e3'�K��J�:tQ�m&"�]N{	��\�7�K�$���xA����Q��Ǧ�	��¾���u&�q��Kpy,�<��bs����v0��E$�ܙ8#��G/Z�u�hk��S�*5����+���[�<+�d�a��|�.m�b����ږ�+��W;uuQ�8|���l\�ʘrF�m�w����Fo�5=9�2����k�vl�6H���4�����t�c���֕5��Z����I��j��D@ʯ�!�zN����(�Ș��m���
K@��`&,��a��z���nr�����7��z�"Bw���=j�b��'I�@=K�2ne~����r68��|�q�v��S�����Qi�p�儝�1Z����P��P��{��t��/�uW4�'J� ����O�%��)�A+�J}��#pӈ���H��7��<y񥂉uu`��V.$-�(	1FyJ�ОO��(z������0�@���� ��%Ub������"4�����uN`�?߿�Wm������Lv5d�Pߢ�f�	��0��5�ب�ם��K<Y��a$ƠՂ��h�.N<li�k��\�)�e����Y:WY�}����Q'�d*㎣��*Zl;D�G�l�	���qW�ج�E�|p������e^Ÿ"1z�	�@�B�v%p^fgvܳU�MKe���Z5���ރ�w��Ȏ_#�2��q�UQ� ���2�|8BHEl�['��1�rq�W��U��td����=9��d��H�3E)��JE�CO+���Ʇ�i.���f����@��}6YS�}��Kq}`\�d�3Ѫ>�{$1$@w×�����AtR�T/>�N���B2/t_� =��J^�;�w�:�������N�oT���s�'�	0���L{M9�q���(�x����^�G��l!���V$���6L���+�E �&*4��8A߯z�\	-~"�˾`ޯ�;���6�32U�-��ذ�*�]��<)f���oH&%����7@��9�\�c>Q��0�Ao�O�c�05 S B���t�;^�0<�%� ��y74��mz@���|d=��%�2����J�`�l�e�P�|ի�Nj�(9��(��U�k�7�vV��[�S]�[t�q�x�y@��u��2��b�\	LA�ܲ�F+ݼ�;����;�p�|�]�;#o�w��~ ȸ߱��v�dc����J�B�� k���Uu�/��wB�T�I��n#	��cz��s���)7�D�������Ac���a*P+�[?7;�'&v�fC0z�/�ʱ�D���}�2�5�s�����E��▧ܿ������,�a:G�V8���6zsS���r�b��U޲9�gm�^q* ��{�#���nF;Rx	��iF��Ҏ|���J\7=��_�т��Y�<��kL^�$~�9M�B>�Q+�qT�j�Z�[{UR�-%C�/x��Y��; �-��8�低�]Q�� �+�_�C�u7��z������v����ƉQ�a.Q�Gw�)�g]�)���r�N�~��+� i�|Q bhѹ;i�T/h�-7��_EH�
Qs
���>N���\ph��N��Gbg+�%���ص
�&�z�t�))���BzM V�'z�M�}-��5�=V^(���t����?�� ?m�m(�{��Ft���tLƿ�k �WF�j�����ww����u��	(��?C&�?A�m�rd  �=�F��Dn�w!(�_�r�vo�L~1�����$/2W6����~�'��*�:IA��)EI�)�N *N"�H-�4^�[����kS�Ci�m�{tN��b	D~L$� ���]$�H�=���ɑSӛ��u'ܰ2I*�ƺ��_]�����G��,лx0uLW�B�����I�2�Ы���޲u�0K�t|� �������9�+�/�S㢶��I��WDh���VY}K&�V)�ˇXi��q�����H��{F��	��as)�r�h
f1!N(����F�pֲ#��P�`�a������*�!R�3�F��S�a45����4:�{`D���]����˚=��J���[ �'�;O��^vS��L��[Im.�)�x#T.9��1 >_Y?neg Ӫ��t�痩�_>�a���*da�+��~�P���r�E��:���q(sҕ����ЈtaZ��%-��n��V�5�`_�������d����<��v�w}�=$oP8�1�ʏ���M8�����u�r.����?���i}�R�7�(75��p!f�Ը�s����1�7�� �v��$ɿ ��Ԛع�g���;[��Z�
���j��jL�F`���d]�jP~lUA�Z�v�4R���|c�+V�H�fC%]P��eM��h���A':��̕�{�N
�>��"���j5*��R}i�m�ƍ$zp%LG���n坵�`uEx���*9���(����d{�xH7"k����D%jO�!�8��ZA���7�R��Uu�Q4iX��Ŀ��M;_��B�L�} ��{(HM��׆��hNJeȟ���HU2�a�OL�����&�'Ciyʕ/�J!9�d��7�U둹��Oj����c����Rk�"l�~�K%bGo�I�*����d����\�Z�h��$�������|#4C�TG�蜫�.��V��m��,�Dj!�E',_+O#T�
f
X��·�[����`D�8�!����g��5�I�:4���7�����K�	�w�<c�6�6�W9t�3r@-V+'�$��;"�^2���7�4{��="�A�{�I�;����4O.�H��D;���2�3��xQ*Up��B���"��`>�� Zi	u���Pb�g|)�ڭ�4	�>ݥԑ+�\o��?=3���ӑ���0d� /�X�SE"E�D�l��Mg�ǉ����.���+cb?���)�Cϡ�ZGL�!�""�#��t�e����q������.3r�k�(?=Ε�B��э2���-{A�����jR��z�k"�y��Xڮ����i�ڳ~���Y�[|-�o�ω��^�*"e)	���gXW�U�<�m),��j,䠛�� �J� �ɀf#'��������������RFb�T��#���9��34�������O�����%�Z5�n6P�ݝ���_���D.���'�-�?ȅ��Xe6��,�VNm�bX��h���8���X�ښ����羡p�?�B�"���ʎ+� �29-���%٥����0��(~Ќ��/�<�4�\[�n ���8�I�r�ҹ)'#2m��%�@����keZeoI BJ��������4�R*x�����@�8�C���M�����O+�c�'��GڼR[��MI _�򐳵5��3x�t�����<uW��,�)�ܰǤ�1DA$�V��*O�Q�w�DhSF�����d�=��g�����M���c�f���!�DA��M��P�b��C���	^�H@����^�Lm��]�y'}<"�G����_������T���>���1L���d�[L���� �P���H�	��
�^�Uy�`�z�(��G�f�����X�@y�8Fǘ/��ȏ$p�U�F���਀���IK�$�i��vP?��ۮs겨7KᕑX�̦D����_N�2��r6>��Ä��E�xā�RCˤ]o4
X�T���<'��/�V���5n��01(��N��
�&��7�gX�_y�!nf�%xH�T�񧪚��A��Ҷ��v�XQ��������dC�o�^<S�񝚒���{ɴ�/��NMn}�K�ώ��&O�+ǆ3�E�nCn�c�����4��r3%��Eb)��N승��f�5��Zle���6�����C��N��k��r�	���LEn��b�"P�v�$���ӿ���ׅ�q%��heE�*%��(��ӣ�,v3W�N���SM/X��\�_�	ȹ���5�G�i����o]u"#c��gYn4�\��	���o��B(��L���*�:�"6���(F`��K�&�Ǘ=�G�ܧ͆_,�LN�������-F#�"�!�^��[1�1ի��-�bsP��p�xi=�c��S���nx7���|T����~�xP�܏M����&b��4�bPMзj)U�q˰�s�@\86��k�$�R�
g.�����WƵ�yJ��:�L8��^������y��3����Ԡ4ޙ��=������h�fuZ�P��LyM�A��}�T܃x;�B ~�0Mó,����*l�%�Yv1��-"i�]ދ�����6���Xl�&ly�^k��o�F���0c\J��Q���e��Gˁ����$)���u7�$�	�6����!� ������Ы���a�E��)�Px�ӡ��k�A���*�'��:�$8߸!x��2�Ϝ�5"KչjS%f�+c!29��-�߮(�@unix̸/i�0?��0��ϛBg����9opx�F��r.��T6���ٽ|#���Jd��v��PK�VP��(��橄�`
Hx	ٖ��q�&H��ݯ�l��i�|I1�� o��J�)��&�����].�� )eclh�Y�C
�^͢�`9N�X~�٭�4��?CF�W�*l)�I�o-t����(��C�z��k�]�xgm'w말%�*��u�6��m���e�%'쉃�#H�G���F���dC_�"7u�R�gQݠ١�3��6P��r�3����,
�!�����bI7>-���a�a2��NkΥ{S5�X�G�bPKkw�+G�����M�j@LW͎&$�g��Z�S��K�����j-�Z~'�U���n��9/cV_��ϖ�	YV�W=���� *����S�G1Ą2Jv��hP[-~}/E�RI���ׇ����Zd���^�0�F�:~<�xxk�d"�B�G�̶)qb��w`��+��{���Us�Y�	uI�9~��-C75'�����֞�����x�\�ڐ+�B�dƣ�5�_�'E-ʝ���
,�����O:Uǎ�[<�l��F6b'5\aK��D�e�����K�\��a\�r"V�@���yd����t�5w��]�+�������ʀo۸ ��_N����q�s[�7�,�xg�<h.���<��h%�!��4ǉej��S���}�4M��"�u~�������u\`�~G��;$֚���Sy�7�6�R��%?_�!���i��дV�	`jp�|;���?�z�(�X6�FbN{ ��_[�=8����0���s�/yh���_���o���a���̌�`� {��&��"�M�\���ܙ��6o���-�ה|�������.g�$���h�� �JG�o>�e��>&X?૙U�w�˛~��C�G�;݅>��K���5� �K>�Y�	W�'�G��V����#���4\������n	z�W�1��v�|j��W�.;��TW�76<�:�b-k��e��Uޞ�Gڱ���|�2f��u>!��#+�L.5��/A؆�����j�,�z���P}�햛Z��fF_O����>W�o�O�@�d�SD�2�������(@�E�헹A������+<�k�I����Ժ�RNv�W���8�U�XT}�/��8A7U) }h����r�. �;+�0ed'���u��Ӎ��<�}�r�]hL=���f�ʻ`�%Nwh˰<9��\�[8���+5� �.u�`�B�:ː�!As��x��0N�)�k��9�]|����K��Q����&=̯�ZB9�X�F:n�8u�#	�w���@�f�-a���:�[�ez����i�O�^���Ꝙ�R�W{{͇5��&���p�ެ$��@/;��mx��UP����mI"-H��������QA~�����!�mg�7-��4��5�K}Q��[i~�<�O1��'�Q��2X�֡K-4P�U�%�����x7���ܾXI�V3�[�vA�#�QχҘb?
oer�����O�Ôr,2��{�s��$}2o'��eנ���d���YD�W�0�{��s=�qb�����U~20X�ecј�ҼZ�,y��v] �JM&0)B0�$-�%��3�cY��?��ߕ�h�Q��-L+3\��*4�:��YS%��+�;Nl��0�8�!�ǥ��*�钛�<�,�n��܄5��m��]��#�4�	6�K30���8zܔ5�z��)�YV�;�2�ڈ�)+�#��M�xC���G�Ls�3-�	(�$���8�l�l�\�cˣ�����qn�
��Ż�y���VZ���:��5�^4v�6������c꥽L-EW��|�LF�zx-p+���)��r)C�϶���B�|opf��qHz��GG��?4���k�T���y�P{y�(8����]ҙ`��y���u���s�T%4���^3_�;"Q=�\*��B��T����(��(�D���L�:[�b��IIS�ɮf���S�t���1�=��|B��\�,� �ޡ�ҵ�WI�c�	߃Ł�����)h�������6f�t��'��#'�����
��A`�J��r#i���:������ѣ{���ӱb:�<9�xB����e��T�����qb��Ν��47fl\�u'�0��c��'o��#.���yA��;<oٖp��n{px���s��F���L�}� .
)�/�+�sHH/N�V�����A�l �����{���w�
�޲��m����h�Z^$ꍲ���m�����fHM8��51�Վ�����)�3��ʾ't�J�흗���J\���tQ�4E~��h���b�?�����_����:c�헁�R
Ǆ��Ek�hË��\��(7"[B�Q�_q��<�~�t1URј�r�+5�n@:(�6�~[�U _��<�_O����ATJ�]<�pD>���tұ��6��a���رΨG�����x��M�����$�2��[��p1�D��p��d����$�Y�5^��*�� JڀE*H���I�Î	�v�,��[���d�<��yz������m�R���w�%��]+ُ޳tH�.˳�
�Wռp4�Z,�4��He��	����[㈫���&���~��Z �%Y!��,��j�Z�9�ft���c�X��R�hLX���֢Ԏɛ΢S���w,��p�6Ǯ�� �7���Bx�Pd�'��*�(�d-�C#[z&�b���u�<m�&]��n
Q�力X��}���_�d+���콶��1 l�˭����R��W͜��O��9��3��G:���(߶V�Es@ŷ��5�˃P�;�	�(��8��?���AnV�,n����Q!,�| ��!�u	���+��d$-� &W���kz�vUW�Q�s�0���t� ���mMh=1u�c����|?��I����Y����Y�1t��Qfi�03~��0<'9�zJ׿R}֑@���X����&��9D�%���*WG �e3+�:��!+}��E	�H�UWҫ���{yK�����'����==i�L�eh��"#�z����ϑ3H-�?=�4���O5~IK,=�9���\�7�>�D�i!���HLɦ)%v�1�/|U~}t��iR��x�q=�#�Nd��+H�Z����N�VJ{(
���a�H��Hc�'��� ���C��Ը|�	��IF8�dk�MLB��1�-mJ��j'�8X�H ���|�U]�;ׅJ�M�1jQ:�# ѡ�Ɠr�O$%w������`�@���]囮�Ns��-���u��zJ?��`��z�*�Cq����>tkƧ0WVD$c�IѰ���f�Cs�Yya����h��*]�^�mP��;Q��'����P��fb_�I�; �%�V��|�nkD|g�����Di|��� nq��VМ�olN�q�-`Gw�8`���w��KU��;���8�E;����JJ�]�M��o�^	��c�"��eգ����mkG�=�������Tq��{�;sif?���C�#��(J�@BxDV�<�|bu��e[+C�ox�]@~��O����LyJ��Z���d��$�'�xn*���X��wiPZ9=�M3!�s�.����,�"U����>���g9z�ԑ��B�~������۝ ]���K��LE�>?���}z��#�1�mQ����>��x`9HwO�e��#E� nV�!G|O�|���'��S�|2�6�ʆ�\�y�*(Tzy�Z�i�~3#Uh�����g�-G;!F��$�AήLm�t,V���	��=�0(�ǳo�_S�m�2��b���!?]Xl�r��>v g>�>�ǒ���+�d�+�|L��H��+%�+u:��; �E@���L㋼�&U��	$B�E\��;%�4��qU��D��H.��k���7��"}�nd��y���8ж#�W�A�u�%��Ȥ�"�G��'�����@���d��|`U����C��� 7
�Xy��Fc���(��W7��d��F�2�r7��������DUXDʪ�ƕ��\)��:q�0�u.�'<I=:�s�ߛ�Mp�	mo�"ߣ<,_ٛռ���K��Gs��hO�R���#�s<�t	 �wd"\q����_D5�_��EZ'�����D<��^*���<08��	��^D9�?�zC�h�VS�H|y��2Ha�@�D!�#�mF�r��uT��*qV;p��������Eo�H�����,*iS�5I_(����#�A�U\_�"��\��&���d�^��H���b�)_��(�5�%T�:є\k��b�Op3wd<C��Pi)�E�����fg�n�i�%��F�d�y8�>e0�B�&�� ��|���C*%,9WA
aI���C-R���L�;4����|̋:AC��a[�^���AO��C;U�
�����p��k�8#ߦ�),�Rۜ����T5�'���X�@".y��f0��j��aUtem��H�����թ�CB�9�ӧq����G5�0��>��{�鋼���̞��g�վ�.	����uR(Y[��q�J)��Ki�aɢ2��pn|O}>?���=YQ�T�U�D���<��XR�+��$/�� 7�6��ˣ����p�;�� �*��E�E+���wL�M���<ˌ��g��ЈNQ��b�U
L���N-�L�8�_����n!���a����K���:ńW|�w�X�I�A�1�Dn��3V�V�N!�\�y���,h�7"�Y�~��"[y��JQBL�c�;$�ǚ�9��mg�1�b&��nX_�3x0��� F���n �MI�@*����ݓlä�o���������2���6l��G����c��V�;����?������[/�)�����9�QV]E�,Lg.dҰ4H>ײ�T���O~��/�6����j%B´���h�V�q��rEZ&��rv��6�?���0��@KlԻ�a�B>{��b��;�Ī`��Z1���}��mWF�EJoZ4���i�*y����o��R���@+��C��S��E�'�S�uR�oJ��lw��Aٲ���[��)�N|#dx1A�R�lL@��,�܆�!�t\!T�����E![,Il���Qa�쟿�o������A�4���&���
NF�"�[]ϑ�Y��v�/��46���Frc_�S;1mħ�m�fn#�h���!�����Hpص��rڝ$�S�&AӁ	���q%@o��6�^�����)���c܃�1R���v_&���%��We��x����k�_�貆s�J{��ҟ��~��3�1�B��,�2'�d�/QhZHP-N���/)܎�sa���(gg�xB^ifP�k�T5��p ��~�t�|��^D|�9,�oo	�Y�)|�k3�
y�>iTȀD{`c��[u�/��K��=���Ve���i�k�Y8��T�]f����N�j��2<��Z�}D���{yvٻ�0|�eK��Y��S̛k�q���u��ǮUK��T~^��7Ql΋Xܞ����I
C��1�TVP����d�v,�vG�����S��F�ݡ/.3��
��?�5OG�hl����������N	ug�J��+V��a!F��\#d����w�;5���Ѯ��j-�����nN��ST�ՐY���k���vy�Ⱎ�yk��ju�n@��f��$mv���e_�����2/�l�=���`D�>+��(���O�h�q��{��.S<��r�^O�Fy�� Fk��d:~} 8�"��wQ��ˏ��:�6��e{����OޯL�]�oe���[�#^���i`+��!��������O�6��|R�rY�\P��x?~ !P.�]gBᲴklT�x0� ܮ��]�ª��K-�[�np���Q+ފeMqV����NX9b|r���a<S�sϴ�J0�`�ܟ�e��)4�jz�f[j�`�L�X�&|�+�������Ç����f���볳��Q���o߄�ׇ���%��댂�d}c:�8AO1{��`��Z;�Q�&L��z&-<����b��?�VP�6�,`�d=�堃Ƴ���������wLVɇS)�,�;�q{�W����0|�G�i�@��=�x���ɶ������$��>�Or�J�Z��Wʍ'��x�C'�G�.�gϧ���������ӳ���h(�
5�f�˼�VH���b䁳E����׏�'��x3������M#^/٘��_@'��ƪk�������2�#��<��f��%��y�c����8�>/R��$e�V��6�����ё{j����B_PC��b��ז�vH�:��MU��I�ю���%k_�7�����2/����s#Ю`�Egy���5���#����bv~�e-�I̵-�c�"Ns1%?<�q�M�����B,�i|�{Ҍ��?~Hum�Į�y��Ձ
����z���궢�������TB\���2&ˍ���mŮ%q7_��W��_"N��~SZ����Υ�!��b;��RW=c ~���}?uo@�J�E�V`�rʽH{�����͹�g�	�a�U�g΃z���7{��˲�n��}�m%�Я8�
��Z�/߸i(�9�I�N]Sl�T�^��zҙ;(��?v� ��������p����lٿ��:eX�����Y�LmA������`��5�3����+3rZ�`��+Ə��Ƒ��ꘝ�&Ҕ .�3'���(9�s���� v�K�ǁ%$<p3��7U�@�^���� ْw�7���'6ޙrQ1�ķZ�����R��bx��I�.��r���J�2?谧$������~�o�| ��,�1J�.�5*�����FD���&K}K3Aߊ:O	�L	E�
�ځL.����]H�M��=M��(u#�M�*����Պ���ؖm����N���������ѭ�v,y9��HT^nU��^Ӌ@X��u��z���ܩ����i���[�!�4��邁�����F�h��P귺���R:]T�X��+4��0�@&�"��A4�p�,�BV�C�b��l�1�Sl�,�ē�u9��އ;�����*�/p���_��URv�!E_z��4R/���t+���ʉ����wfb�~	�PeJ��Bp)Y'�v��b`�łM�m����!h.�Kq�� Њ3pFV�����N���+�Ɍ���Z��F��AG^��-�t��>����:�wW������&cO�zb�cJ�=�1�Z�S��Uò��D�BQUK�%�_��.]H�$�0�׹�9M>���>��#6I�4P�=eb�g��ky��K���s�����j�d8�aYH{�D��/q�D5o�P�u�3���(���^�{��3/l)�˝�����3O�3���f.c�k��Hm�hS{j��f6h^�����H�U��O9��by쩄���;���-�����~c�.�8�((eE#\�-�V�:	���z%�Ǹ������ �d��a�t~�������;Q���fM{�����Fq��	Ҋ#�ĸmV�a"��$������7T$�
�/��;� ��s�B~$W�	��7<�zz�����c���(���Sw[��e[L�
�m�k86��!��[u8���T*5K�ڃ�%u�E���}b阰G|��m�mۙ�I�!�O��FEm��j�aEt�����}f`�����*h�h�T��13�� n5L�p)��&�!oy�˦���Mj�����_�y��y�"�%,�"q~���)%IAU&�}ί��?�S�m�/*��4Ja.穋G^^rO���<�g�QO�F�5Ѵ%��ubs�~ B)�^ɐ븗(�l(�Ǩ�\*�&J��8��N��k	sn�|N�e���n���[%AZ;��>�jĻ�=j�ԥ�~�GK,�U_��� k����0��Ox^��M`���`UK�fqb�M`LiX�� ′��p��/�׵�fN%řڞ��0��utl�[�=���� �d����<7���z⛃�Vj!�J\�e���ɹ�r1:)�l�on"�8K��뼤;�	D�x��Kz�u��~���ĠM��5֍��%u���g�Mr�JJK$�b^c>AZ�UKM���7��Q��6��/�<>���0��EbKp��ܛryi�JU��k2���KN�6������C����J��s>�=����~�GQ��5p1 M�m�n)R7ǃ1��)!�Ĵ�} �������`7R8=p/b�T�]b�ܲê�Ԃ������д�XƝ�X-�ǧ��5�dhĪm:���i-y�������>|Q�ml�?2M�!���{����s=D|���^�b	��Pb�B6�)��+	��1e���?��	��4��(�a�/��?�q�o21�[,��Q�$�y՚+��9&����;��P��L�D��@���ԓ��v�����I2��b�B���|��0�q�@�y�H�1E�]c��H�خ]����^�����8��)�����F�[�xq�Y�Ӕ2�w�D�o�*5K��\ڤl�����
H�]����J��x�;}��ͱ�f-��4��M�-���K5��v����M��@�ɹz��@�l��;_:m�2|$���x���a��h��\�&��*|�VLC��s��ɶ�
KN7wC!5�|Eb����yn�N�ٜ�E3z�����	���K��R�Bwe[wQ��^(�c�8�P+I��dӜ;:����n���YY/��t��X��s�9N>�x��=AKi�2"n��:�U����%`|�:i��[�pW�D�� ���5��<�t���Y1���HH������Q'��Q�
`���r��s�JZwo\��"��i���w��z�aek�N}3Ko��u~��[��U����O�mUg��Z�����~Ip����M�{���Y0����L�K�c}g���%]r�cTB�7��9�u��ۧɔ���
*AbI��.�-lݚ?Z��+Zҽ6�p������\aT�Tʖ{����k_��]�/�=�Ɖ�����C����܈)L�XSɰ��"`���.t��o
f�@Ju�����{���A�tȼ��<�(b�>7љSFg�c�x#��*xyT��0����ȵqH�b~Ǎ�J�2;j�����c��K�J&��\}𮲸ivʹ�pC0��kژzF����2AVNmft���$)��C v2��q���m�H����`Q�$��X���H6ݹF*(�ښ���)�ھ$4$�h�s�{���p _�����l��U/�CnoHP3k *�_�Ǜ_O֢��w���<؃�3nWs-����׎��5${�	�W�>	P�%.3�v�ܰ��O�vG����{�ϦR���h���C�[�f@�pQң�SǍ&#E� &�|B�F\������ef �����d��G�[�Lq��Q�ZiV
78���3��x1R\r���t�*�N�1`�Cl�&.��L�`�V<���P*�ǀѕ���˅�>���eQ2?�`�@���'��'����\��Ʋ�������	�P�v�Q�h�r�٨��P_z���_��X�o��R/�w\��5�o2�?5|4�*1�Â+��� �B��D "\����C�F�
���	��I_�v,�a*�g��)��~ѥ��]-�N�E}��|�~z+�4Ib�:D���1ԯ"򖼲�Ն�����͐�����h����F��L/kь��z��i�rX�]����/��7��2۷������-��!;�w�.u���G���H1��O7�EX�% ��cvi��2���U���-�V�s�s^"��E�"�b�d@�)94V���Z���%�o\#ד��q� 9�:�����U��u����_5�^f�tjO�#��N���>�5v2L�2mI��B}�����S<�;����w��<��/���C0e4a�Y�	�=��l�ԧFvo]`J��.��>�qUǍBg��O��^�.�^���\tyj`�(�dG7[�L�@�(��`F^�������Q5L��S��!���mM)�Y��!�Xp�bA��ڗ��͝6Ѵ�qp�E�Ӣ_�\ٮT���2&ļL��	R���DBA��
�#�F76�s\q�R��q�gdU&�qap(����M-�ꂼ3m�A�%GB�BЉ��o���C	>��̵�˥�l��ab?cE��b���HH���<g��jM�)��
�z.p��z�3k�w�1 ��g�b��� ��KJ�g�9�w��m���e���^Iߩ�!]J�-h�	c���$��L���+�	ݿ�1�~ҷ?հ��yT�o��Dԗ(c�}�m�7}%=ߧ2ye�a�t��l�3����nO;�B�	���5>zF�*{lm���i�����M��������B��|ˉ�e�	؄�^��@�vV��"A�+��괤s��gf�}�?������. ���v;yip邜θ�'8=j�����7EGHFk@����a��V��L�&10�2V����$'�hC�a�2�M��
�L�Dp!%��4���=Pl����~������g����هˍ񣌑K�>�o}ۃ�ܜR𰠧�c��o���O�,��絬�0:N�P��z����O��4B��	+g�����16�կ.�{Xv���kC�1/���輐Z�9��i�Ğ4W��������R�����׆���-�tGܫ�<9�l*���s
T-��.1�V3��f�i�8%a91|�צZ:�ơ&���C�J���"�Yg؍�C:�>����'�/�w 	�1��d�l�f[�t528ڽVj������n�����a����/�<��$�zQxU�`9C�w��i�q
f�Pc���M�\����&�Bq�j�|�.���+�+:�nz��B�:��ȧ�����k`0/��g�v�����{/��bz�r,���ol��*�b.{\h%+7���Ǹ���ɮ�k#JZv*eD����!�a�"��?TN�1��2*A��12��l̝�6��l|;��!��%>o������Y߱v�u7�B�8����cj�[з{�,�9���gpo2��˗eCD'���{<^ڊ�ʕ'�?�x����^B��`EB�u�Z]U�y$Gk��J!rh��j+G�	_UU�6Z�o6���#�߿C��5��[�r�D\���g�Z�+-b��1_]^��k�2��}�H��9f��1\���}#����"�Ɣ�Z��,b\~h @�����Q=[��j b��_��f=]lB݉f;��>���"��9��$_��.�q����y 
��/�.��3KRڦ��Xh�i�@��)����њ\�8C_��bm�^)P�j����X_nRұ?/��q�����4J��2�/��sI�����2��ٖ�2QO�|�8vNoH��u�ܝ4Hb�9r�CƗ�8h�/�N#�AL�t�.�� �\pѽ.�5�E���n^�W�o���t܈�y������oxO�*�f��pg�b`�}�o�7|O��'�~	��dǐ�a�˭UݐRp�������K1�?%�.�/q`+��c��U��)�=ՉO���S���\ @z�Iή���
N�F'jPl�	l��a�	���S�k���1�2qu�u�
7��u{v�C3�쵎N�|'�掎J;n*t{��y^]��0|Kdn�:�=ҴH{������~�) �b(
эE#-d�#��]ZE�\c��rt*�gƁ����lT�-��TA�fY��c��6�I����6�娝y����͜��a�0���ȸ�h(2�D�\�A���.bx^��/T�n��Q�*�[���q�'R�.s�3��u��6���}+X��vކvǭ5������5������̀
q~�ݗH���$�q���t�Z�ӈ��!6��wg(G���F�^`�)9׽gń���+;߮^����2�r��Bvo����*>��ED����Ȭ,����5f�\�j�:jo�O�v����u��V�W�P��j��E~-Vi�^��$�5ĖJ����;r31�az@h���ы�N��\�9�g�N=ÿגsnK"H�=1&o���#�(�&�Wf4ɂ��Dk����5g �u�3~p�g���1�01GwP��!��P�;�b [��3��F
��-)�|���#�{6֗���tM�O��'�I�E��͎f�&��8��;�8����#�n�0M�Ƅ�ֈ2�t���b9����g2�*��5Vp�,|���L�ѓ�E������F��l*l 1V;	b������A��h�/Q����ʯ����⁣�I��oX� �d�m&���b��ӡo���	�3Ȯ�����Ů�N �h�i�>[n���Y߭[��X�I�$Zg�L�]T��E�^j2"
}l�F����W��PY	�:���υ�TV��>o�m�`s:���x��E��ݞ �wl�QB��}ft�����NvFZgtQ����R	͡���>'khܶߋ�������Hyǹ�TK�&�'�q5���[J�X+h���#b���ap�f�w]YMX�v�7e"�4{@T��#��ͼ<����J�W���̕�(�!�H��.#���Tn��f�����ndh��n�/���)`�f;���C�1Z
pwHW߰��҅N��"F��eiVD���4[5���B�@�`²	�T�/��(�F�DRAՈa߸�n���Vk��Y��_Cz�j[SĀ�=Ts[����:8M�R�r��򲝤,*R��(%tH�����v�)�ȿ�j��*qc�@��p��I͎,Ǘ��Π�Q!��ռ�F��1K8e��N4t�-��UÍ��|��n�b@�-�'�x;�Mnd��:m�؊V��s�R�u�T�g���?A@�)���ki>�c�%�(\���E}(�(��e�;S��p���zrpc��~�c����Xe��W��)��
"�����I�|yhz�qh���nz|�Vm�_�M�,^Ɩ��3�T=��+�K*ܧgKӰ88I��F��PJQ����KW|�Z�h��*�����#�zAq�D6V"�����[�E�K�|Q�d��7�
PC��bX8 wV�>�m�s[Be���"��e8d��Eq����/�1K�ly'�����+
񭗟��t�*O6F^�|u�e��!T�5��c��$��#�gs�yW�>�ō:'�yV��G'@��w2�Х�|WY�F�~j����/���߾u4w��X��?#CW��"cb(@��a|��]�������y���ё[�t���Ք�
k󚫡�S��/@�-��a�t
�p̔��K䣬Ga�aH6�t59 	���>A��HȔy|B!�`K?��h3Y��`>߇�uE�~�d�����xh~L�ũХ��0H�fL�P3N��I^��n�C�b��(�q�uX�K\�����:x[$�j*��d^��$���'a��y��r�?G\4D��Ĺ�ޢK�kz�9����Z�O<���+8����L���k��函8���X���eOo~Uj�P���9����D��t�"�=\��/����~��ɑn$E[K1�jn
�c��5���C��3�߹hX�d����i�U|�p�.s���3`l�J��b��5�a�c�ݐ-�@��D& ��{���)��3�(�~e�_c����؊+!�Y��e��T�z��4��Ծ86��{����c��v��gqT�8{)!����2S��8�x6�ecrkm</��~sG��:�ة3�sJ�n��ξ.i�8�'�r��%ln��N�
бr+1V�z�D�gVl;���nb+Z<0��ͅ�a���L�_���P�6��v�X�L���|̺O��M(s�E�a��Ua9�a`��,�����]���~=�2�ђ�d�daC�ERI"�U����@͈�U���ތ���R-M
sp~�-(�>vP� bNK��Ů�%}AtLL�֒4 �rvJ��_�c)���Q�gq�^����ق)���#�����?n��`x'�@="�l!�|��4�ą�9Co;E�����`�"�'͢�U7t��v䳶X��Ju���c���P>�C�Y���4<,Z�Y!�Y�E&�]x,t��B�����)E.i��<7 )�U�j�Z=�VAV�U&Y���@�j�Oi�����6�]{j��<�73���2��歷�^�ioT+���dn�tN^])��r�k���SS�6����b[��a��[��ǮgZI��t�}ͯI��UY�ω�7�kmhF߯م g�ݺ|ϯ�jy��%����S\� y���Xg��S�ށ5�<dRyEu�a���P%h!hs��_}��ڤ ��OX����;P=��F���� 1lx�
����W�MO�J0D�!�W���Ϧ�\�����U��|(��br)�G>O�@IBb�Q��QSu��K���|AU���Hz)���JlZ\O�K��gv�m=��EN˨��J��Ӥ=����Q�K�꽉��`�����(���J~Z:q
<���Z	�A��Kz��Ǎ�|�0�<:"6F������_�H��]X����ʸ�h&�
���J`��gU)�q[�c�F�UV�iI;��K��q�N̔�j1.[*�z��1��^9�ڮ�y\��*$�-��BjH�\��&{�IK��;�?�	w�����U�W42��?[�q8��(�`�m;�<��.P��x�+x�\�8�!�q��l�x�{�v!��M�����<ժ�p��g!��;t���q�wJ-��i�?؄4�)�4Oǉ��!*[�O�a��r�`+kiS3Nц �����<����,�c��͖�FUl.��ͼ����^�q��������	-V�e�H��� ��`���J��~`��H%�7l��A�{-(vB_�>�Ʋ�H���˲�SB�'[U˒�L?��*h�|cj������ ��P7�RmI�����G����~u���Ё�Wܛ��p-z��p	ڛ�}�n�q���*
zfe33�00w�M���8W+V�(r��K�P�:���ԍVN��JCp&�v9��b���Z���:�ɚv��I�a��������L'����3�;�:�Ƣ���Ti�`#T�w�^�<(_���(R��a�2l@��s�U`��n��U�¥�r�M��'~P�&6�vf=�ʿ��K�f�������f�H�+���2���A'_��=��G�j���f�7*����i�,�c6�4jp@��f#�"]����ӶQ�v'(�#\�� H��]��%2�eߴ8�2L7"[?�;�HF��j���ρ��d��""Ȍ�t	�Io֞��D=�͌R+hID�.�&�p�?H���������RJ��TГwm�X�M�t-	���b_0c����#t]�6(��`jDLE��TQ�C�I�Gq���tU>�$�lY���Jk���$B����'��kg�,�Ƥu�JBJ��+���bx�r�������{�L�(�)j��m�*(�V-��o���Uz%|�.[坡�iM�O"��W>�݂|�F���n�����a�A7::'u!��G�DK���k�0�2ʀ%/�h����V�j�΍A�^]kx����w��0)�'S�:�S��\<��|�����]?j�_X7��\3c]'#�H���GFF�i�i���RF���ߐm^Z�%\e���bt������.�)Bw|�> ma����������� �����{]���;��1�=�N��|���g���Tk��E�~3C��%dI��U���] U8�ә���IS���1��u��[Ut�_�V좥sC�{���Q6S�m����X�P�#{�i�:��;s���C3��P����\�GA]1>m(��x���3��DW&��������0��I��E��4%0S-G	�w�̡�M�z��\�A��+�m�˾�U�¨�B�˘Ю�"����6���eƣ�J�ὦ��u��"4eh�G�j�U8��������O�� �n�s�V�)v�{3�7H{Ɋ�(`xIdGIT��K�T1�eR_H��I�T����2�<ܯ��2����3'�d[�8B���%��lv/��q�VN�{��64r�S/�}��O�;Fc�P���7�c��&�N{����M����%u�!E��[��?^j�?��qZ��!���޺��rN���\䐙,���Y�������b�A4���@�8_˦��*�+����f)��,#�IpJ���74zX��Q�XtoFx+�C�an�j�g�`�8�h��k�b�w�V�-)ē�B�p�$��)Yc�s0S�.HO�5��%��.����e"<y��JUIm��9GR���j�&�3/�֢�[������g> kŠ�4�ο+o�ʀCm7�Tɐ�8����.��!���8F�����_��xS��j9�|ɴ�xb���bu�P��.�_=F;ܔ�6a
��TxNJ�	8��������8��E5(����ZF'W�57�2��.��H�z)h5�D�.��]�	%� �M�z��g�.0&�:�=���l �������y�=�#P�<�5��K*C��-0����K��w*TO.�U����0O�?+��^L|"�	]9ة9��㕙���~Q�%8��rG�Ч�ݯh�`' ���_�����(��M�0�T���'��LÓ�C^]�{�btq�QjlT�~���XR+wG#�h�_�{a�HFf�A�0��ڻg�9p���U���^�_�r���ʄ��U�AMާl	a��8�}bV	�ǯ@�'�2Ym�$�a3�G�-	�7N�����U*���y/�$�:�Y�g�7��T�#�d�{�
|*gcG ��l��4�����~|v��.���Ke>Gir�����ē�P�Šb�o�o�i�;az�p��O#�##���~vnC��!����M�M�%�&޿�Ԡz�އ�#�Ķ
���]Y�POC�|����G8�HyX�s,� ����@�h�������u��H�/����!�aV���H��'4
�XX�r�c���N͡��M�S�0?QW�K�.�9Y<鼜����c�*�r(�8?���0�ŋ�W�O�~'�Z�׸hvv�ܺL�����b�7�\+�g��78��/q0��]M��OYa�����t�`AL���a�/�.;+�.��M�۵z/�� �VO<�Bx6��J����}��A��o�xN8�!D��׀g�#�>d�'fɠ���']퓊D�W?HL�}��@!
�cx,��*�����{�ć�����6MH�ie6-v��(&�W��(M?�����8�}��	�j@�[Lp� �VH3��:�sq �i�:��?/���Q���X�A��L��K9ưgl���wf]>�F��h��Mp�P��X�u1�<��ف��=�V����pf,�Mb`:���R�I�&?̛V�]����M���� ��.�,�|�U��fT��͞U׆���1����� y�g�2;���HnQ�G�^l����B~��].#���Nv�|)b���g���c�Ȱ�1ꪖ�_"V����.���'n�Y*m�^��t��j�{Qz�=?η�<5x��v����"(�n	�lnΰ�����ɴ߽�T�l���BYѡ��v���iO�~ZEQ��""�&].�� �&E�|N� ������Xr��j} ���t΃_w�d�eJ0�Z6"� B�;(Z��N�(��5\���
�z�`�� Xƀ���0���B⟐ �#J{�&��:��R�1�l,��_Y�"g����F�VҜ.;�F�?ڱ]u|���'͆�5N<v�x����� &�]E�"�+�|�?�z�)�#(����+�C��~�9�W�͵�y��
�K@��(���b�Ur,�X�Z�j�xn~`T#��̅��L�w�u�{�i�Gt�	��J5��Y��z��'�Y{S�'�����ta��9enJL7Yc���Y��3�E �򅲇�;�Y� <2w�,�$�`*eWx���E�EJ*�{E�S�i�`fӈk�GLW�9�LGèض�Q�$��ͣb(�<�RN�S�nJr?z��$ΰ�����Z�5�]�;5jb�p���;���Lb�����uք4����0�ˢ�Q��+Ȟ<�A��NY�=|�R�8�c_��ɣ��H����¾�>��� �ׂ�����۱�u���s!�.B�A�kP�4��]�R�H_a�wE
.8�ш��)���劺�k�L}�W7���Q{ٜ�b���Y
a��Ж�����i�q�Ďw�^�ն����tk�Q�h!�هh1�Г��C���g*$٧bK�q&	���L���{f��]*DӢg?��A��V�LdU���_��b��9���qЅvk!�ML��v�؍z\:	��{�Ei��Ęs��bQ�=�]�7k����aM����[��j��긤��^����2����)��',lÚ4�X�) ?J՝|g#�eq�'�,߳k@���έfS�o�w��<�)�����X ���n_B#
uF������2jd_�W��*jQl�✽��h|���4;kf��x��QR���Q��E7[��H��=炙.���Q�ڈwK�@�e�����pq��t�e~g$�O����Ð쫐�Ŏ~�eK_����O�Q��d;ȵ�S��S|7<w���~dܡ����p����F�a+���F�%˛����=�	�B!-� 󲎊����F����S�����ltA�"���`�!�G�9i�g��F1�@�-�̋�ۓ�N	�E�a2u�[;(q����q��V�g\�5/��*����'󄰭���0�k���7L��/E�!��-���لW�kr��- 8�R̐-,Y
w(U�aEݤ��� )�6��!2����o��0*�⇺�fA�|g��lx�Kw��ɗ_*	+Z٦ac63Iy���}��_.�ZT'5�o���S�S\�Es+n?�t���ȹ �n�E*��S�;�Jq�{��I�A���������Z�����{H�ʪy��fi��fy	��D�VF�O�}��+�X�^����Pi���ٌ�_�^1�q�!�etM
��'Kv��w�֮��o+�
�U94}��#��-X4����Х�%�`�͘�Y����Q�I�I��W/?tejM&� pF��:�h%����)����j�u^ݣ��븐fz�۾ȥU{��ދ�YCnˌz�z3"��l��ʕ�<,N���>���S�E���("n���u*@��5��{UwW'K�Q��(�����BJ�5�<S..k��i�or�=�����b"����xhNs�����CJ�=���-Mp��I�-{�G�Ҋ	h�Z8�������"�:k��'!�%�A=n�	?T\�+�]x|g��F���>W�;�@�:����i��U������� �󬂘���Z�dj:�O�`_�Ja��SBK�>H��J$	�*�ϥ�tl�b�����䥵r ���`8�;����.��깆4|;J���r����"��(��,ۥ�͝W?0�zsӼM�N'ڹaj�����n�=����3}w=�#5�2��=���9^��	�X}��^�j��2E���N�r�ҥ^ ���)�6F~��
3!��� ��;�>h� ��bb��eK�������9ه,)f|���e���X:a~���]cI����9��{�������"�N(ׇb��5��:��i�	��MJ��nv��6M�D����O�57,���a����5�a̓��O��+ �n������@ޡ�R占ؼxE�L�*[eF��qhc�D�WXN�p�b߈}�6{<$f��m��v�T��N�d�$\�,��ETV*�	��ϑ�S-ײ5��*��&�Et���Ï�(���=�C0ƿ�`Z��~B�C����5��0�D�?ag�I5j��+<�kծD�B�����Ae3�E���`�	�HWj�p������L��*)Y&
�8�b�A��)^ԭ��P?P�,�)Di�>V�;�7���VV�z�~��`>��Oϯ9��i��z����%�Č[�T��t���u �O��o��R�6Q�6L�T
��H>Wē����h:Udf���~�(%���Z ��I�����:��	I��\�D�~���g?/ӗ�n�B��x�&��|����/ $ưU���)�<��c&��秄|�/:��O�Zi���9z߻qp2q�s���&�._ҩ�_G�ޏ�[�����G��X��
���N@K�����T���'�3EV9cR�1�e�9$�,8�+k�0Iݶ"F��N&��Ѐh�v��p��5�ٿ�w	���k.tH��
�x��k���_Q�"n�X�	���ww�~l�\���5�<SLt��m�\l��W
k�!(�
��g���1�:���O�K�3��nNK;DB�[郱���6,~�.��{�L3B)"�_*����6���uq��#�e�/-�l;��zn�k�v��Y���j!e+����8��Y0��|مm�V[�.&��n�ր��se�������dp��%Dp�Yt��[���� j8��m^�[������Ǖ�O��݉�kt��(����|��a�#L��>
�4j%��%��Ƚ�
ճmm�Ϟƕ�^ŅD�1-k�{�Dn�!d�g��W����y?��)[m��Y��K�k"���?1̉��zbeB�ݗe�`�N��xWGhf����F���,����o|�h��,��̐����d��7-�Q�44�׉1����ؔE�= .*�L�N�����x&z�AOI�_���VO���M�=�L�W�J��l �O�E�o�u�Xbo�����J�c�dQ�x��4���'p��k3��O%pT��rP�[x+/�l<�Zy���,���ٶ@��\�%$��w(ADm+�,�����Y�[d�mg���x<�8WE!��2�Td����#��F��℮�:8�e�'�H���Hv�{�M:N�\`�ڨ����݃Υ�j�V�L�����ϖ���a/��@s_c3�r<'UU�����djEc'n��E���)Y�2m^��h����m�
YIN4
�bF���k7;�1=:4tJU�[5�:cVV�eB�%��-�"= �z'�u��z�����İ��[9nJSp!�c_>a�Ryeg�5i�Rq��-��4�Z#c�0��n���-w��u���)sה��Ӵ'�>�٢υ�Lr���փ��x�I�&���*sm���S�J�7�c ���N2�gQ�v���<�"]���#�c�N4t.�'����8���/ �^O0��4�5�v�pS���_����8��
=�ꇥH�\H�6�{�CP79<��Y�m��G ��W@��X�mP@���6���f�7�2��ٴ�8��	�!3���A�T���|� ��g�Γ/�*�" �	sU�=䐭��fqY�0Ld~z��ހ	𨋉�oK��� ��ri���M�<�n'�ٮn��S�>=b�Ð��r�������)�LA����ź�o��ۧ�f��2gRz�+�;���'�1�H�7͹���+e��I �E�m�B��-��6G���	��=����8�yp��1D�w���ʹ�P�F��T�!�	��l<�>�01������xy�7���a'DZ̥��R��hn�����ZxP�~��6��/� �Wq���ɦ�ai�HX�0� �=y�Y/+�8�Nx�ĭ#����-����U��0S�g)�i�S�C�T�`ת�L���h�%r���n�^w5_t���b��E-㺊�Zֶ�Aff��?<@�����ޯ��5�uU��nOԦ+4��90��|�H����@���}X8S���������^����"+���ˠ/�t�	�:M�04�X���#X�
�ܾ�(�c��e��`�u�TfN`�;\����JP�v��qF�_(b�����+w�+�-ys�keu��º�~.�b!�v����`�G%dOO��*���!��8d#��lմ��~�՗UT'M�<�WA�����;��ȃ�e�wd�fOMӑڰ��N���!�E㠚o�st�g���j� �|h}d��5�)�d�Z/h��_��]������}?��>]OQM�K��t�T�|o[���RZ�T������G��Q��I�'�� s���<��6�B�p���Y��)�<��h ���?�����\7��ya���Y�����oxp�]Y���� ��2:����m�p��sz@��krz�v�gI�E����L�d��6á�iX��o�/?��֗����v~U�2����lL���P��\�ם��9�\������pk	��S�=�t�4�HE� $�	��>/�JA�=PN���|Qhg�1������6�2X�OeV�0,��BSV��%#]�pik"��:B�����Xǆr�d*F�E�11��:��"k�b�n�7�ø�3�n��~ *�!�ޘ���-~H�DR���/�f���m�nЈ<j��Z��MR�w9��V�Y�C�	D�v�#�.��|z]M���[2(V�-� �Zj������d=0R�	E ����Qk/����OH�y��>��V8�7u�iB�i{#��KA/����@��:�X�5id�h����ܨ�){M]� ��2K���L4Z�����]T���#���`��Z'��:I��0�Lf�CB�X���[�Fzo�.	����}B$���e۫ɔ�yq�1�@����t��.ݡp���Z�����J�h����9rZ����9�<������,.m�-�*�0�-)��+�kS�,G����̍��N7M0�r"C�0��Ma|/ ������l�[ ��7ޤi9=��	�jX���!sBX澹Z��rl������/I�a�œP4�:W@�ҡbR�{���'�Lu�ծ������vs�y��GDgf��+ز�e���_y�Y�ع��Wz������h����_9�]��a��	_�BF`&�.��6fL�|c$�߷s��D�Xf�xKelp�'��2?sy��*zT�蜄N��dr0�5�QЁ��y�����ݖǽoA7CgX�m�p��;��q��Z�f>�~���y*�Զ�F�X����>7���0#ޝ���`�[Mp8�dylq]x��p���A\0I��-���h��i�8 7��W��W��@��c`ӗwb�dotM���f�?�#�q��Q#��t��0�6e�cx����ް�]n5��.��*	?���w���"����d�%�L�dCO�Z"	�l;������]2�By����"�[�s�ɓ�ό��9 s%�
�!���Q�<%,q�4��G(�����vYz�<�ǸN���-��G��梭]u�X���+ּO���?��w�:���P&F����g��#m�{I7�f�_�% >��J�ZB�Y�$U5�2p���s�EB���z!�}�ľ[*�B-�'0�)��/R��j�{۩Zd9ΊXR��d�AT[���w���W��̞�?`���@����_H
)��dZ�˩e�6�5�I`|W�&�.�h�-�� ��VW�������
���s?/M*u�[���}$E�HM �孹��̣���~h���ۅg�q�J�E��1��93nn�H��0��q}+�k�7�l�.̡�"���z0,}���L��1�N�+�%��������n�-��2���`�
;]]T�A���cLWߨ1��7���X��I�5_�80����<�{w�ve4�� (D�����l{LSOGc�M��������Aa{���]%�f�K].�	O
���?�ȏv��mD#؁�u����rI�b���㱶��\p��H #~���i���4�O �#�1V�l,��T5���=��'�@9�$�i��G��GF��H���$\��a7Õ�B��=�Y�l� c�1p�Q|>��S����-̏b�;-�	�w{w���S�]3�C�k��@8U����uI�c�2�4�v+���1پ����_���W�g�EOrC�y�h[�����ƻ��g<�\���܍�B�!���}��-��Y�l@f�|@?���
Y��&
F��	�}������h��u8YY�m��6�����z���pl�E�(Ҡu5T1w�'H��F���"��>�h5�ps=�E� @o�~�'{����N�-&�*䣥4�Fp�ET��~iC�yI���}W��r(��E�WP�D5�+�O#mn�䱘��	�l?�Ҥ_�M�z���N2u�O�(���t�V%����u���̦�di���_"'H��[���G�R��1����ɻ?�XOKF{zd���O�y�U�&d-&��O���S �)ޘ����u��G�d0E���怏k����5�������/����ր�h�׉���'3ʮZ���5�]�fWc�AcX'�����n��͇H&*ԛ5��;HGc]�B:ձjh�`���(�F�@���7(��<�� N���� 
$��V�ݭbO_�.D)�5l��d���w~���F{�E��WiQ;�����Lh�ب�޵aʰC�½���9L�ͬ����@�:v�^�õf�a"��d%z6c04И�k����N�����4�yzp<��&�~a�����.n~�UK\.�F51���_�E^��P/d�g��F�X�� m�H��|+z�|Ƌv�h���4�)�2Fx�.u��s�7�}>Ph��B�хK�bhz�8��AgĴ!J�*ͩ	��gx��"%���J$�	�uO�����`�3��Rd�����}�Ӧ�	�,r:\��[�&���+#U��i�B��yr�ͦ��g]}������	�Ze)�6�?��e���s�t���(�����Saz�J��ȍ#��by}�����^]}��P���'y�YݰFGڟNr|�h�'qND(1kL����.�'~�`j�gd�$�j�l�+ԧv�Zͱ
��5h�G���v�E9ha�r�c��9����cӠ�p��A1� ��6���ٛ���!uq�:�#�~	�
Ϩ�G�GE���}<ǉZf���Ĵpd�J
g�r,8���bҘw%w�qg��'�{��V�Hf ��C3��;<��F�!Hc�m��0�5���D�/�AGo�N�=,�R�"��w��pH(�9��mnYw��NN�8~�&�Ŧ����Wg+d�u�_��Q2S9b��"�C_Q��rӤRr�8U�9�����s�Uڀ�{.{S�/o��iɑX�S��!�<d��li�3�2G+ש�ĝ��@�gnM�JzI��ػOW�2P���Z([Oh��_��,�z�&�r���ּ��=�Յi��}~�Ar2�Fpm��^�MXyƋ$�H�#a3�
��i��Λ<\w��	^�e��1;`-w�.�'ܴ�;9���ǡٵ����)3����~)���B�Q
�ȖOˏL�u�̤��!�VM��ܡi����f4����h���B�z��4��b�<"v���,����{��D��U��	{Tz��7�c�7K���`1I1�\���-�� ��u������X�똬�����������#V�Y� s�lz#-�+ƅ��{[P�yp�Ka�i�V=��k�e��b��R���L3�3ӛ5�s�V�*x�퉬���gS�`�ՊRM�5i�d��SWȒu�7[������W/��n�9*�?Y�����~Yi��
������/r�Ұ}��o��������%����JM�����
�]�N���ZDFZ�T���z��S:��[�ys�~�X1Y�����e�)]E�� �_@���k�m!�N�)*�V�5nty0�$�{��(��XV���/eVB���r'*�6Gu��f��A��v����ܽ��gc;`-��\u��4���(��fv��(Q��������a$�^J��4�����4>o�}0߰
�y˰��/�ݸ��c��NFh���?Z1���8:�HAU�iGY���$��K�k���Q;�L�gI.�X��#O~��p�(��í5�j3�=�se3%�c|뀀��AϟW��޷\@�}��!="o��oh
�j�RA��
�q��!y'��^�3	�p̆垴�E���B_M���;�H�����bW�R�Ἠ��
��}�)���,@
��DwїI�A�x-ݔĬ�ڵ�RB����(m��?�U}X)�A���n����Zpy�mhm�!`�O��߬��Q�m�E�3ƫ3Z��m݊�e�B%��j�"