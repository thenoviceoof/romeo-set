��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�ϗ7�#���H�����u�g[iˬ���t|�3���ҥ�ys�B�@Yq�"F}�\"QY����#�ڇ7�\ӷ��繟��1W�k���q�u ���{�m)RM�S|@�����ͣz��yʿG��O�Yg>�s$h_!��-~���=wx�=�M�����/�mb�K#�� ��1��W�i�{,?�EM�N�0�K
䧣�:39ok^�(��-���V�f���Sk�	����}ؖŸ�*����~������6l@ޱ����t����_.��±7�Eۨ[�ܐb\T�8�����"��!'���^C�he�K�Zw��J�;��E���a�BnB��lje8�i�U��^w�K�@ܚ��^<'�������������a}��a��W��S��!�P�:�ޓ��|=ǎO�k�σf&�_ K(yǦ�+F{v5�X�x!}e�y�D��"љn3]��6:�Ѳ=&:_��h�,�klf�es�4�=|��-�#3��r�E8m>�e7�{�~w���O3��{	 X�n���7��[��{d�mҫFG�6�ݝZ���4́���GF��yw�D��Օ��挹O����[�K6���L���ڹ�\Z'�
���lS}d}��w7�� ^$�j_��묡X<P�`��&X���xRq�y��G���R��B�}[�b50t��j�k\��Ju�a�V�ؒ���w�\%RF�Z�購�:*EO�GT+���,��B�/�9K�5J���t	���y"q��yǕR�<�]���>{�t�f�'z�(*��l�����'J|N�]�F����Yz�ȅy��/��)�B��
�vu`o9M5|�Z�e������gM"���C�W��f,�o�`��<��Xk�:�s#�T��/q�PC���k�!}5������j��b%׊a1-�b��\%猢��S������Ew�Z���UYwds�i��;�IT'q��z9}j��!/m�n��4�Z������ء�\��0d��>�fZ{�>�Q���}o�x�/=̪Y�I�s<T�y-���G���_�җ���2���5�g�$K�+�'y��wj�%��� ����s�ٸe�p{��V�$C����FQTX5��)w�"��c��Lg+Z�fvV@4�ZP�>l���
�U��������tAĪj�k��V����>lv�C�/8��M�jR0�:q����Tԅg%�L�:�����t}W�/vF�XȰu���*_=�Ҧ�/W �W�J��k2|�v����Q�o�2�l� �@��n�S&E����q;�Ǹ�(�b�?��&�pAM�� k;Eb���7��U�U�k�и}8�+9$��'����ݧa#{�~P�C@�u`�#����]�S�N{"C=l
�i��+*<�L�n�k��STA��s�%�X;�y��@����L����n��e���-�4���=���t�X�	���B�`�K�C���Ɍb��8!5te���i� �������9�E�y�w��ܺZz�
�5�_�w�.W%x���|�	
�Z�� /��x���f�-H>��|�)O�(�x��:E��&��Ͳ�Q����<>�E������B����
\�t΍��9��Ȟ��\���$�z`�� �1n@4/��e�P��$���u-��?�J�$?���Q�Mʕ��[��y��ن@0ha,��t�H���OD0�p�{O��M=f~-�G����(*��!m�Es'�#�A~�G���yk"�ї�����!A.���Qձ�&Yeis?ޖ`r4��9��7H�͚J9i�Ň�yʣ]��,�y��)�Wz1����?����Wt����� ���� �mT��"�\<��o�����D���^ϝe�x鞾�F̂���ˁ��ͪ΢:yz���Jc
��CN�!=�,�]$a�����Ù���2���rTc���Z�=HZ�$�Z��^T�{)�ȧ���_ׇ߹k ݧ �dظ�z����*����D��٥=ɬWb�	օ�����^���Ar�pLPH�7��G(�.O�]\��Snf�ǯy��(za:e�^������.�Ƭ�r}�GMP�s �Ǭ�����O�x����Y�T��3��`��3h�s:����\2�d�;n-�q8���FW��>3�|o�
|�ÿ��F4I����[Lb�8��9'�Yj�l���[T��i�V��p���eƤ��h�9���`=����[Pf��c���#����4�7����Y.@�ݧ��{��Q�MDm��D������C��2��]�4���vK��B����s�6'.s;�Z�U�e9J�:9�7��@T�_��ꐜ�M�x��>�`�� ���"�k�(V�я�����5��GS����ׂk�M���I	ǳS��Q�N��P�ĜF�GA���Wy�j-���D�k�*��M����ՒJ	�q���Y۩>q�S���R�(Em�F��\���-�h���Pj	M4oı����DN�����(,�,�|��SO!A�5��.��2�ɉz�	�K���q�'�=[ʭ|LX��Q�h;vn�S;̝�Є�%/o�f?*���[�B*�z��K4��)�D�gz��+.ݕ��c��%�V{X,,7+M�0cc��;L�W���zo��ϖQ���"�L7�k��1�鲾ě@�uo#]��` �00�v�3)��e�o�g9Д�(�e�$��5�z�m�7*'��
�.�J��ly�L:,ۨWu0B٤����?��RĘB+%yY�|�Q@������¯C>�<卓���<X�dI���I:�!�r�4+#(lpؒ&1���эb_�+V"������a!!�h4�B��PS@ {4�i.����eG�\�w9v��<��pp풥�OYY�0������Co�gFFp�[�|o�s��u��-W/�Hx�o3p�+F�;Lг6]6b��$�^W(�,ބ$���(�?�g&kyt_�e���s5���VE����{l8ݎ��Z�x�'8�^+��Wl8˧N�]v�Xѡ�t �m\K ���a����)\�$J{�[�=�4��h�}�iy2Z��TDy2@��k�N0��~���qt�x)�{��N<��LW`��uT�*���(�;�)��)���@N{��'zoT)G� B|e�eH\�(8���@�,�V�6����r��_8K�E:��&w �aeC�&f.f\*������2�e��C����<���
0�?��u\kYA^M��*��i^�X	��0]Zs��))�z	��l��8k�aNe2��i��3V5��]��zv��� f�\��$��Oƺ����Ni.�q-�Ӭ#��X�	O6�<�)��c�Xͱ�3��X�Qw���8RJ�x�(��xsC�-�
;Տ����px��'lHR
��Z��{|�{�1,
 �e7ų��	f��������~�GPV�S5U��0���(�ẗx4��������W��H;�*����j�;��������f�������D�Q�H�Nڡ��gT�Aw75��7�:�C�X��4�>�<%�i�Z;n5�VJU}!�0��zu3���ky��`0��M��
��j����eqw��T�xvB�c�1EzhMP]0X�X
"4p@HHW$�ik\9��D�{����i��Ԉ<�2M�v���,�@-q�%v2���,�=��埱�lѕ#��
%Z˓u��O�
�q�:0m����K�Pu�!0�;���j�\�Kyv�k[�0z�GN����ժ��R�Y8-&����i�]d���� ǹҷ��c�&�qO�&o.F�Eg�=A#%0`�Jn��U5�I!�d�l�J�J���V2Ylie�K��:_BĘ���;�����.B�|d��`�g�- {�y�Jl��L��&r�6 x�M"�p{�[�{Wc�=�!�ٓ.ۓۋ_��I[n^�� L^�
��2���I�R@쒬���H�n}��ఉ�y�fÅ	���>�,r�-�-^�<1�L��$��h˰���L��X�ibI/�K�J��jXc�n��w<�A�J��ȅ?����N�ݤ�z��5H���ߺ�=x��S�ˉVH�x���Ր����p��O(#	�ӽݸ�� '���⩊<0�v�o����V*��Kr-�I
�w		Ŗ��i��|����9|��N�3�
(=��0Sh�@˔��f��Un�6�V5Վx����o��B<�99?P.��/ H����gY#0�<	��� ��+PZ�E�V��)�J
��s���.�N�ΙyŽV���_I��O,��`�'��<|��YЗ�[�QҨZe�T��B�0\�R�:�&�>�B�Nݠ�,ʝ����/��� u�=A����#��d�
z�U�x�5����T��4�sK���m��E5�rfcg9bx���ʶN��V!�Y������)#-D�+)��9D�$���+iV�9�SaP�	�p�~>r�o���n17�7RRZA77e�)*D���˄ߣ�d�f��������)�%��< J�v��)4nO�D�Q�)�wDX5�@a��=�;�7��a_w�OR�zw�r睟�;1�?���17�0F4OaQ���܎��Fk��bp�k��o{��u�������?z��dl�+�H[m��5��xg�#3&4}����J4�
(U��Q�-���3x�T&4H��(����|"��Z.��
���hN���Llk~n�q�A��1��x��Gޓ����bt$���pԸ�P��K4Ķp����w�Kf,8{k�dA�i�p7��֩�i�~}�G�d�Jn/��1?>�n,�i~�n�sh��D���g)O5X��u$+�f���V�z���\(xL՝\�GaIrE/`;�&���m.�7
�\��y4�Ie^S��/u���V1���?���B�e[ '��{��SB� *6���k��� KR����z�����h��g�x�ǭ�ʧ�Č����J;)s'W=w���z�9Ich)=�_�#8�{���\����=�/�`/����ԂapQ�����X�+�^j���`0H�t^͋�Z���u�R�Nl)$�^�w�*<�xG����.����Y���Qp�wu�y`����R�Zj��@�ery���y��	ܠ���w���$�]u`1�f���pd]ӏj��u��&�fU��¤��7��K�>^FA@gp�
��J��N�l��[P��k�Q�����Fy���Un#g	��g��'�mO*��P���N���1�>W��c��l����Nֈ�=��k���6�fsm;�\o��m$hjAW~$��a��o��`�@�c�=7»9u�{^��%�ؤv�F|{c�;ǉ+ac B�f�R�3�g�S��J�Z8�)р���F�OA'y�[��⫖%
�L �0�}żА�f���,^���kи�>l���Hf����j��G%�=�ܣr����dYD}q �y��Hf�
x����F���8#�B�R����s�[�m�Ow�C��"���F)�ޜ6iP��k��ӹ�z����T�;�o�Q���×HE���n� ���z�f��?:N�s��(�j��W*s��u�f8}�U�K5�#a�5+��V�bKI�R�K�rQ�a|�U]��xq�����n���]&%�\�/�a^�:�3Jkc�'l�n��ǎ�5(0Hש-�u��J�z{���@�1Wӆ�̀��������VCQ	K%kl�b.�<�Sx����c�Ü�B�w�1ڙb;u��Ʊ�������50X�hr2�G:�����JI�'�IO�V;Q)+�V���.��wh��.4*�gH:	�(7-��[X�DT�L���j,ӏ[���e8�'xd�O���*���Yrnx(������x&,K�<���d�SU�ߗ��J	�7��J?H�ڒ�@�f�p�"ћT�#%�E/}�K����>:E�����k�R.��Q/��7���%�ʪ�b��|�/1�b���谕�TS���~���*�5GKf�/qk����F��TkF'��ReY�KmVv/����-B2 �`��j$����M�FGC�`Y����EB�I�e����P]N/:��9�_�����N.��s��s���4]�aI�5�
�l��N�M��5����W�!�]f[���h1Ħ	��Ń�_ZX�l�է賁�U^Y�E2|��lƉ��^[)�G�����8�%2�0X�D�t��¿?B�O�7���ū̠�8�N�"8�;-�j!����Wk�}/����ȳr�6�(�e�}T��2�U�P+@ސ�ӆ���AϮ�R7D�D�/+��oC�1�U�#�i��_p�4�3��G%�]#��NwN�zY��Vۧth���������TL�`�3g�;�e�a�@L?���t�mOWX�p�s:�V����a�����C�!_�I�w�)���a�������xُ�+����R ��(T�ierUc�4���t+!��cO0=n��+�CDp�!}g0��I���jH �A;:.4bYv��#�w�O���c9�@	�K�5���Z��
�$.��c�+���cr�3d��$Ч��ˬ$�G�-��n�%L������Fdi2������t�H�y�,���v �$�=Ͻ���9��[��r��5��9�J>��T,��X����ʟ��EQ��)|,��C�]8�����y|dާ*��D~����#Un+~.�$�x#b��v4����v�=�Ohيr_���1敾W�	������p��1�t�.4æ�e4~��"8/V������|*������贼�((@��]{Z��H�� ���\�s�w�G���q't����[!`t,wNV�8㾽�-_q3��hD�6H���%fv-��4���a8��5�N:�)�[���_l��F�yXX�������+��x&`,��Z�`��7?g�/b�ɀ �9����/���o.1Ʒv4k=��z����Xn���0�Y�4!���A�!���mK�{��FE��Ww8��qeVd(�%J¹���0��ܹ��;L#0ݱ=���]P�j��"]��i�CC�&�GZ�VY�+#C�a�@E@���2�� -"'�xf��s��6�mY2.	��P/�G��$s|��AU.�M=��+p«3TF�Y�@t,�Qb
��5�Xj|�*8��n4�]��ii�l��Y6,c��1\���&�����k���e1�m�<������T�=:�#��Uy:2�� a�C6�0�gܛ�q,Ix����Z����-�e�JB� jnJ`��~�1�q��ڀ���2�j�Q:�@?b��1��;��,x&b '�8?�`S#��B����&��iB�]@�L�#�/o[�oI�
�:�4��o�ͬ)�K���@��
Nf<$���m/!�"�׏��3� �����T��Ƒ��=��y�-�r�1! ��1ix_����v�3BR7���I�]��)PS�ҧ��f_kA����Q?m�������hc���P�z%��,~k���w�Ͷ��Ξa�Q��ܪr/�t�EuP���6�f�������a�����W_�J@KL�9�`�#��-疩/bl�FW!1�����*�����wZ�)��f���ԃ��J�A�.�h�@C'�����*�T�~��"=��rL' �vC���I�{�- ���&!K(�.�s�����P-��4�Fo���E��w�s� ⢽]���-\O'�߹d�U�	�jH��ԝf4�;rG*D�_6������~P!Z?�;wА�T�T8]�_�>�)M�����tXz=�{���4��rץ(i]�v��Lhϟ�fś!Y�K��m#�/���~�J�	����*�o#\�H�!>3}-����Nl��M�m�__o�`���R�5���R�e���'5Q�Yo����Ø��ԡH��U��t2�o�	�		�*��c�lxe �WEmK��z2��347Ԛi���䩰��bl�Y~��f��Wؾs�ڝ�&Ϳ�	���~'k�gC'���&7K� ���œ9!�;�Ш�"�9����SrEƷ�������Wo0�f%l"�A�M������Nx�9�~#�-Oy�e������Yʛ�=P�[\�o���)ga.�� C��߶gk	w\���w9~l��z5Y�ڻ(�`��,�U����<����kd<"�Fk����i 2�*߻�����m�i����*`��Zɕ��:+�5R/�,M�lb�O��.�� �s��ۓ�e���sY�j�w�P�ku�bm�D|�G'���I�;{���n��&�&��{��4fk+�[���0#��u��%�YǷ���D���ޜꤲ\yjK��~Ɯ��1l���
������i49��\odf��'����$�ۤH;�R���}	]G���T��uZZ�{@ߒOzQ�TY����!�z����ī�jL�n��m����4�sEu�Q�-�	�,5ёZ��C�*uɇ��?'�G�;Ek���ʣ�[��f�;l*�д�#�斡�{��߂��=���"�z��KR��r8]��D7X(�ﴥ��"K��$��|Ao&��v�����75jV,Nh\dΞ�� �I�%h-��C���Yy�1q*j���qN��~������]gG�L�m"k>�����:\���٦' �O\����E���׊���;��;^&ժ�k�P@�·3�z�eȲ-�N \�|�}"�h�e0�����'M�`�x�R�U�"��6�ܳ��ou�ȋ%C��������I�<R��������N�@��J�ٶ�٬�u>;����x��ýCۦ�25�N�S6� �dS�b�y������c���U>Y[|����W�D�;c)f���YY��ELtN]�wg]���.T�c }�f��$tեn�����Y?W�NO��8�w+~]_�*���2�x�e�bq���F��	��bp�$��=5-譖I-3��Bj�?"!�v���A�Q��	��%��c{>o��!�Vޤ����j����b`�P�w}� �dJs)׍Ci�Ej��$��wk���\�
����.8ɲTݑ�^�h��L��?�F��a.dZZ�d�f'gF�7d^ h�ۈ0�I�汓�=�|��^kla+�O���N
�+�S�>zxM��d��U�P��{C�L�Bv�v4̿����q���\��k�G\)/ Q砷D�ǌ}��I���1�&�����ZtN�*�H>d	�3l�V�@��`]����Q��YU��1�#K��?N&�=5��|��ž�%1&���u�)�T�ڞ��p}8��o�����y#�)�����5�5:�'�ũQי&�'��5h��{ֈ��|Q��8
�i �'Om��CK�w��=Vlos�n���a4H&+ؕ�n�{g�|VW�W���LÌ\�Ne%΄�X��h/b-�k	�joz�.�Sn�k��!Ƭ��6���Z����5�;��x@�~Q�˙�ɿ%��='�3�{#���{jᚱ���r�f`��_��+5�&Q����� +M�/���g�@�񡰧�Q�̽U��ꜿC���;��T]�a%S����y�e�e����5:	����b�m�.��Z�5�;;�a��EZE�o�N� iީt�������V^7d�pr���Rʉ5�R����W�5C	�R�y�y<(�wH�o?����.�Qp�DK�}&HG��38\h��/o�\��w<h���Dd;_�cїlX��D�^$/�ۭ̐ߠ��E��?��j�Yz��OE¡՟!U��@S}�G4zj�m=tr��0����ۼ H
�hՄ�OZM��B+���S�(��<��E��>�J�5D�k�0otN�T��Q��Gh�6���^ѷ����3��p#j/�O���� 7���n؈QXܢ���w�u��c�AX�^O~��'^�I3h]�����4sώL!Vr�7��	�g<8a���$i;�
�{0�p*�}�vv��#q�9y}֎6b���l'�Ә�D�Y�EfX�@������5p�����s~�������c�?�4��Y����?��*�s�PK2 �x���x���w��)���X��\��f��K��""�Cx���y�$~�BRvݧY������*�xUhnrY*��Z�U!�%X{�
��T�F�H^툉��s�
ncX�춼�7��\��w�v��$�T�)��w����yp����ICXuu��H�f�:�ִ���<�*Ӭ����9���
���B�ž _�ݥ����HH(C^�#-;��KZ�%�ǐ�D>���?���-9�9<Ԥ��u����_��E�[ꇘa5/Ia�f ����"z^��}H�`첒-�k�)�u:٬9�8U�6�ݎ�~A�E���D��z�h���S��b�W���A��n����*A�%�sf^ �2+�{�by��uַ�#xt�~���*� eT����N�d�����ms��+c���
[�*q�s�*��d,�b�M����͕��7�h���e���{=#�����]��0�I�q8n��h<�P����Q�O���,@4/lS�PZ�ar�&����ƕ�X�=��-P<����&�c^��d��;�`��Ve�^�5����'"'؅�X)(S&�z���J��<�vT��`�'�q�Q�a��%��6Ϳx0��hȡ�pO *u�-��Q��	?C����u����E�C���O{R>�;�Vo��]�J�~��5�:f~. ��r��ͥ|s��9T#A�g����.�����~r������96�7SROT��R��g ��KԞw���G7ߣ�6�u�tn:&��6��|l����K"�(�&�|� K�'���{|f���-ؚWy!��8��?۹�K�\�U���b	��v
�l�������WWh���x�H�����es��b���#!{%����*�-}�{NwK��RۿiX/�Z͜p1�o��nma��-0���;+��t�a�j��4Մ��i4�i��X�rp"���W����S��d椗���%�?�g/�9�c�p��x�4�w
�7@Gpr�P������o��epvRK���J��Ҥ?r����''x+s	|m��;�v���> ���IYH겆���6k���L�O���3 �^a�%y��P��+;��u��yg�`��+k\�������p�=*y�j��r�
��C#�<�^r����V�dv�r��X����!����сj-�[���.�./��T���;^����/A���0�r����3����q#��e+��V��E�L��~� ��h���}��H�]{&k>*��l0�Ne#�b�)�ҕ�8	A]�{썌��*�ʠ<�.K�fVe�fS��*63�5Ӟy�4��?�R�9ǟj�1��_���Cb ���PF4��@T8�e�����1߲H��W��gY{���)�����і+ח�lgk2�������6wq���)��v.����Y��Q� �>	�&q�`�����S������g�e��&����&6^ོ���ir�.(����r6uJbF��\oGo�
�bE1P��/�;M��6-a|�A��T�('Q!
�T�v-�S!�̈́_�9��b9->oM|c"�Y\Tn����df��+�*����-�:ni��jM�7座_��B�^�u"ͩ ��%4�s�I�s�z������z��c[�4��˦��7����+�`���S���#g�~�`�@:�s1�g2�p���[���k�$�V�ɲ+x<h&�#��fp2�A�A�7]����Y�W/%G�I�1W
��\�s.�Tu�t~kdW��~�-����Mh����=ܟl��QV�51�SX�,�]�fHWU9�h���oa�՚ ���
J��t�!�;H��~}i7�<�t�0c%D�>��q&;x�F�d�f�n�
�w�Iȯ��i7D�R� 3�p&�%��F�m>�E+n��FI�eϒ��GT�8F]?�e���rV�"�6I�W'ĉ�&dMP�B�5���5��:~��A�=j�2F�(Ø-�կ�?�|e�#2��W�nE���I���C���Q,�oe�շ�)b�!B^�h�km���L���(>���Nk��ۉ�b�Z�/e�TE2�Ͳe��6`dv8��k�����Q��j��Ks�E��q�W�Uc�"�XYz�w%%#쬏6Tx�����
���L�� $��>�;�ѻ�������ϧoe*���S�"�ǩ�E��y�8$
P7!,�E�����
�!+�Q9�c�*�@o�D�L�߫Q�Es�M���<�n��7�F�t��A0kI�Pg5����0!ͦp~i1�lՉ��C� !w< �� �}�����o���v�ҏC(;������`4wϪ^��An��m0�� �=?:1���e�-�9�mՄ�CL��g�e9�>Bv/82,�xgS	���@ ��Ly�,�����;�L'bzϦn!�g�wG^�f,c�N�/��	��N<@�k�.s�\���B�~�7�)c�GM6J�qW�]j޽�Y��Vn�ږη=yL����o�]�S6ĺX��c/a���(��.�t]т�_P�G�<c]��/�L� ?�����"���N�upwMٔ+	��fD��N��e�L˥m.��`�9Z�۰C42�_
J��B/��v�XU��L����^r�uv�r֪�-Z��v4����)r�ۣ�:4�����?\��eD�6"�4�̠-�����!V�Ug��y�9r�ujpXϽ��a�sP.h�JS��T�]��B��v�r�.ѕ?��m�'O��j�S9̌v���4������6�X�8׌��H�"p6yYF�q<�����Oׄ+��nZo��h�!�[.��b�E����`E��K6��n(N�n튱���2�P���c�'��������V n�
�]>�e��˓����O���fP�nN�Vgc���w���h�QBm�W�N��T�Z�wCX�����W�#I��W�Z�i���^�,.W��(A�C�*A�,#�>aϵa!�L>ۅG;f�=+*(����]����ϫRV�Ƭ�Ǟq{�gY�������<! d���+3�>��[�)m?��N��z�QLZ[[(M��w�ʱ�\�6�b"�޹|1Ȼ���FV���T�DID�p$+aoc�P:�t͉n�����a� 2�G�ż�����O9�=��I���T�1�S�Žp���rZ�0Q��NK7�2���N��vD�ێ�z��$2z�T�F�b��@�@o�;�I]��y���=�3�_������yd~;"�<����Y��P z�b��8Y��l7>���ϧ{�(+�q�Y/~Xt����$�.��{Ǌ۲F��m�4%Ѯ�����*	@U�"���?j֞Y�+V;|��VH���T���d*���S~k����_>��������#e�	wC_1�&�ў�!���~͹���[�k��2h��{h�UwW�>|:0�nȈ�FGe͒�%��'�����e|����b�]F7�Np,r����5Fd�!2|?�����`�i>VMT��X1)E�������p�c��*��\rfݽ�c�QsmY��J6	�q�׋V�fK%r���h��ћ���ޣI;�b@A�S+�Rqb����o_"C�������W�J�/����59t��Gd������b�<&�9�ߤ�$�N��5Z}�����U���W1�ӽ.~�3
?t"���H����T�s|��Y6�d�����N�q���bN����D��ŖL%��b���>�T�ٽ�4%<C�>W��f��`s#^���@I��dl-|�׼��0��&��K=*�G�C�kX��T2�k�RMI��Z|�����ݍ�j����6T3�����^f�p� ����~�U���:7;�f�S'ep��^�N�D�Bs�����k��%d�laB��O���*�����x㚶�wbj~�G7a���� ��)I�?,?3р�%U(M���%��6��!$e�"�:sUX;^2=�x�h��frș�����>	e�~]�U�1���\�:�2R���A;]�%�*o��:���N��Zy�T�����`�=?���Sq��JW�O		{�- w/#�S�H�P��/C����?R3|���й�zmO[똿dkfS�!�޳<g�V�a����t�N�V-� �eȪX%b�(�)#DoN}T�xNW��52Ӭ�܉�J�-���3��'���r]�DyGC&�����n��Hk�9O�[��#�����̣�%�w�C�+x�pi>S�ȑ����������~�'��+��Cv�m��IX�)n��R�"����Ƶ�S���)]G����[����IF��Ѿ
L̺�Ke�J��,�i�APV������K����a����D}h����S0EAKTCK�]��j��?�sd��A<C	åCW���NE��6	aΛ���./>��k񊯚p���&�?G�sO!,>W{��v��w=��ZJSz!*3��1*��Q���҃�0�ڐQ��m�Hΐ�3-�Mx��\�G�eQy~��#X�4ϟV��%YH�7a�0�7P�\`Q?��5V<E�*�xН��r�Z��[9nv��Z�Fb���e��8�hd�����+;:P��	�'�O����J/�e����ޮP��w�t>��k��	�����=��ɞ�*��H;`��Ǹ�*J���b�*0ko�7�W0^քىSKVzה+n�����F��tk�wh�e)Δ�m��ʝ
�Vv�k	�����
R�*3\<jm�P �pX�l��m�bڪ��J��^��������6wq��:"�TQ��(k��A�m�VlD�o�7g9�Ri.kD�����Q HdP�/p�Gw�PXTEB�&��/�dGCn�������u
�63��T��� �����{�f !;t���g������R�8�6�a��k����]��ܭѴN2�gt�6A?��YK-�$���@^}<��m9(��#�����cy!$o5:DC�ev�B����F0�'�s�1HG�	1o���Г�X����r��>��.�IPY���5�� ΃�8�\�A
��0:������_mbE�nM?C�J
����Dm��e7sAs��s�sfR]�!���F/�C�8�ܻ��)ҝ�?�s[C��x��TvBN�+.�J�ǋ��n��nkK;L,,�{L�i�i\}pB�T�B�S�}���-�M�*����0��#:�j˕! @��Me@�	9w3��`�a��ޯ���B#ߴoҵ�b~������Z� F,�ŅҾ��Ē����q��kJ���_�)��Vv�ת?
_t=�2t�1OoH��'(+l��^��`+��7��RΈ�0��7&U�o_?��'?�v�0���\O�!�<raa����n��"�_8�c�Ժ�u%~;��Q���kD��K�%V��E��^��_�W-��:lUđ���3,T{�V�Ou^/YK�x�gD��d��"3�HMkX�?�|��äje�=��;9��;��h#�f4���k�u(e���h����g�ȍ~�����e����᳸�hS�0�L�Ӵ
�R_��PE�b4�C{�99�ky*ɮ3��*���±�K���7�G�dv6��>��ہ�l�'�_cҌ�� 60��ZR�@n�j�m���꼙9+�5�*��E�h�'.�CC�6��f�|1�Ǒسp�oȬOL�N����.%�Fn�j�=cs����[���S܇��S��
��v����|��o:4i�
�X�<g],�{)�G�!��g�uV�3�ѩk���ٍ���D��]j���ғ
xL��;#�i}NxR߳��*5:I�Ȫ���� n1��gy�7��FW�tԩ�AՁ�wh�ěҬ� �"\k��#o��]���"��UP�3a]�,�ү�}@�I��RJ<�#�1����� ����դ�@o1#߻����ܠ�h}�o���3>�r�ks<�G�r��<�@�	#���
�����D�J�򘩴h�6��'��ȏ�sе��_Ri��%c�(��K�O"*AR3ϕ���)1�L z��l��~�Fu?���@Y I��<ʄ�a�'�͐����1@�|;���gw}�����X�7��)��1�9|�u\���-�4�^���	�A��]��m���l\�Nc�A�Ãg���uk��8⿈=��>�� �ܟ!EM���j����K�,��ߕ��"�,4��3�o, 3k���b諽sN�E~$6���>�b{��lɞ�����`��Z,���gB%�&lX���� ���E.��覸�ߘ_�e?&�]�� E�pS�˿Q#䔬���WUX!]�v���LIw&�,�7�u����ͯzU��6��Ȓ�[�'REd�\5Д�dϨH�H��, d7Rf�>�c�7�<o�\$<0ܪ���_9�h�q�IA�Y��*��o�l��eB�M�?̅���c4�D��PE��x�tDA����W��H�[D�ޥ���Q�>����\n8�z�!}���@�#n(�N�N�������\�ך���<���%���3��?m]�QM1bW�����d���xL��vnYs���;�n�:����,�P��TZ�e!��#�;t
��꤭��vf;� �=e+�&N��ߺ��QY�D:��-�p8v|I��N��˭�7i^ݱ>Vf���j���,�E�u��� {�N���pOVb:�2���czhl|��YpE��+�DG�����3��[#����*5�f�'�fl�d��YZ<ȧ�z�͸��q�3k���mg��!��!NC��/��9�����F�>w��Yғ9�={�l��,���Q��Ϛ���wޓҭgDP�����1�����V�1M-0��^�e��/�:�HZ��beQ#�(���ǧ�Π�i���f��垣��	�P{�B���9�('�"O@9qX��7�� �W�,�M� ����g5�I��r��Y������٤x�P�[��
&�h���ә�bU���;���HoHg�į(�W�c�#����`1�{�� �r�̺D#9{��<������"����Z&���r�>	����M<a��}}7xh.C����b[;k���3釮�mԓ��aL҅����ԯ%\������n�9v�F$9�56�n�dY�sq_SCOw�UY��?� ��T>��\����F�����tE�|������a��N}�}i��&3�Oz��AY7A�Ӕ�/���f~�&����2��N-�H;�(��IÙ�!t��Uؓ�{M���hM����e����ʙJ<�m����3;�H��
R�+̇
��??�̵?�ߒ�/��n�:]�9��h�� �O�p�l�V���E��^�]�mʨc#��+1j6p���S�"|G8#jf#�ԄD�R�F��x��d�;�ɭ����v5+�z����Nk���fZ-۶��H�6�O�J����V��[Ja�q��3��e��_�����"� �[�:��|��?D�D�[���=��|��:�0G],�B�t���n��M��v~̮��G`WnHY�i��О'\g?�! )ίR�k |㑶ё�9��<E����?��Or� 0�T~y ���i�Y�R/dy<Z����j�{U`(�W)ǴGv�RW~�ǅ"�Ѣ�*����R�e��n���M���^�Fo\7X����y���KN��Д�Z�
L.�7�a���ڟ4 O��G\
��{��7,�u��	z^S���O��I/�w)[���5�sZR���c�̚�C9ק�ք���ҡI4!��!��D��7�Ɂ����-�2�]䶙��Ə>�~)f���KU����8�[-�ЃY��� ��������$����f�W�8�p���m<_�G�[7�A��P{O.|�~��#��ik�����bʨ��Z��T���N-ՃJ��U���@�CV�-�mP����yU���$���,A�Cl���yd&�'L��=^�Z���ħ�G&.h�	4�ۍ݌{��z��0�f����*գ#	�>��c�sP��
O�s�F�����R�s�����ܡK���b��!��r1�D@�L^ɔ�7k?�#�N-��|܉��]���(ғ42�y�T".�;�"E:���3���܂yŃ�ό�Rۆ��s^�}���3T��
�uG�����_~�p0�n*�ɔ��pl�K�R���`�H �gT�����	@���*E ܇���2��{"s:��~�}V��?6�u�AKW�{@���Xv�7
AivEQ"��B��T������I�I��]'+a	�L#����U3c��Nd�|?Aw*�E_�o��F�A(]7�GY�#��]���U�:�v��.K�d�1�@G�ԥ�9~���H�G����]f�T��r�O�3���O�����%{BU��ղq.�&K	��v3c��\Rw�fH��b�e��Z0v,�l��G cP�K��N���<��:z��
�Fj�!�r�(
��;p�S��D���x����k/��fn��8���5��\��Mv�_e��sF��\SM�r�X���1j�k������*���=�N�,B>�:�5�欏��1��Ep��۠y) [��(�:�O�t X��_z�%;~+
����%�F����y��A__k�cqm#v�c�	C��!�8��}x��ܧ�����%��V����cʲ�y�/�����nGƀ@m&+��ے��7j`���QH~$"�_��UD2m��e(I����"����he/�JC�5ߙ|+��S��L%,Ĳ�	��v���H>H���|I6��|Q�Y�)DTd��ĭ}Y,#~���2�櫣�VXp���U��!%Q�L�\�pa�U�p�#*Ue���sx7���$�C�r8?M��)��X�<�J)]����������\��8ȻBվk� LM�%ߣk��h��Q�i='Q	�b���s����*Wo�R]í�j��܍q�(:�Q�	(���c}��1�*�|�&�A@����T4�i���l�����j>�o��L��|��b�����r��v���� �~}�>��yL��C��SiO"QOӛ����ţ��E`�:��_2�|���k"�+g>W4(-�A��1�%�pM�uן�X
��dC#�ϖ�&�S��0������{���5
���FSE\6pg��Y~ Vxï����Ȭ ��H!��{R�5���]G_����%%7ɯ
���S$�s����/�/ȟXw����P�x����6^R��p�#�g�<��p�fc�]�f3����4x8nW{+ X1�"	��Y-��2]��Pĩ��n�)*�f��@}��;Y"L:��kj0F(�%���Q*��}�Ñt>+L��dw��hB�.�xEH�h��e�D'�CRU$�p:�^I� ʑS�7������%C�@e�LطS3�f�Q-�ρ!��!��#C �o&�R�=������r��5k��^��?H�ȝ)�$0���o� �(���J1���N&��� �`.���H,�~����q
�K�S=��FW6F+�C`T�$t���	!`�0��@�\���$�,���:;D,&;�@,��!h���ޕb0<lO�7�s�����T����zx��{��C��z�I����%䤇1Ek�1��aw�SWm�|�S���Iv?�����
)����7Kα���و���=�
��k�#T����e(iR|_9��P�Ng�.��+:��g/-����u�;�'C���=�[����k�Ơ��S�S�'����[��K�CxB�G�TX�K���³̭�`:�V,���^��*d-Y�yD�s7����l@ �#�m4V���9�{铌�]����j�o����u7�I/��4�q�*5��b���r�k�i��L�����ܔ�WV�l�J��Ƚg�\\�'Hn��Ѫ8-�]�����5^��o������.x�*���0�zof��6�XoQ��U��f������6� [8J���9"v���lCe����A�97Ɲ�и�u���I<=��	�G��O��f��'���)�ٯb�R�SO3;���ެs��KE���oW���v��p�.�J\W��m���h�N�� 9X�71g�d@"��<\+�=(�2�}���~�|#ub+!�i��_t�������K�2�>.pu�C�L�*�w���"b�>�M=�0:��3��3��4HdU�!?x������X�G�oR�zҳ0���5Ĥ�P���#R�q��
9��������#i���l#]�� �NM���
ڦ?#j�>�	��'�= (��*�6����;�D��!�����:U�Q�ZGm���c؜JTm&h`��м1����y�69���&ȜV�a�ʨ�`@�V��{	}wD���6��.1�;W^Z���l���-�����"w p��d��4�3��P�߅e�x'���q��[�
<WAy�5x}�]oVf� �_$W�=^G�"�6C���������<O�| �\�8%������0�|�9 ����	�I��E���+�9(�
� `���i�XB�B��cb�[���HX����<�]�� J�zYr��6^��UX�ށ9�G��j�Ke)���eŊ0VA���&X�
R�I��,X�Ϭ&���iK��o���S��� $!�o�'�͠X~�͎m�����&=��P�2�ۙ̓�ݔ�t������ﭦ���{���a:����N�]�m�Գw��~�������{��i��6}����񛕎��	 ��1Rf��Sgyb*?"��]�k#6�Ɩ���m8��O�b��T�����Y�L��)���~�vu���Y�7��CByO����9420�Ϙ[��ߩ����ռG=���Ϲ��Ph��3Uz�'���̪���`(N����'��:����DJٝ�k0��ju�����RP
u�����Ԛ��|��7=zCJ�c���eOb=	�.����U��������ϡ|�7,�Ss��Ss���#�7���������kL�;B[���2՝�0V�m�\8x��\���J�E�l��i����$0HLCt,��#[�YvE�.�!f�J���]��H���m��D���ٌ�v��&���d6�P��>����Z3%(�2��ܢ���}@�q1@I	�QnW���A���6�4+����d���T[[ycJ2�z�-�W�V�� NU�jL�&Է���l���j+i�#��)Sa��_��m�N���]���7��=6-P0-�@<��a�z��3�݋�D�]t�S^?ye:�/�V�������Vt�d�ݥ�E{�����"�-�ηsqw��t�W����'��D���7�Ή��@u��*߅t�Q}],��qB����#��߭*7��J^YR\ů���,7���@(E��8k&\m�+�؃�^�f�5�2��G
���i�v���}�}f��hR#��i�	�Q��n(��l��կY�*�e��Rn״�u]*P�l��i]�G@_�K�3fR�
$wd�j�.�vAXi ���v�L�_��p(�t�=��1`/$�@�?���<'�Pv��~����.4�'\R6����-�s�S�I2�����k������M�5f�Zk9����2E�hra��G�� ��O�M��Λg�	�@m�t�9B��� ~Y��r������� ��;�w���٭M2�M^��� ���B//	����1s�&qc��ͩAG�23���R��W�����蓓�;�yh� �9r��l���o���͊��.M2�̴���j��ͧ�^����<i_=��Yў������t*͐�Jp顝��Qم���~���;��o����r4AL���&�� � ��K�R'���d[]�x�dtw�2��Q礑��t,�v�<�e�=��r�O�)T��Ҹ-�F�׺i��Z}5ݿ����/l�)d�(t���ߨzWh_���B�g4�k@����9m1�Pն��"�^����͸��P�9w��`�&��^�>�Y4Y�����3~Rz��_?:"�O,<;F���ʵ��=*5� w�P��+Q6�g.�tZ��>F>*��-��RoJ��3��
�w`�
ty�c���:T�4y�{ϼ�$��fNrc����]���(o�(˚ �!ls��aW�A�����o*���0���ǘ4v��e*)z�f�p` �R�Jp��Wi�����D���GV{����2�#e~�Xz�yo��K���	��V���>�?������"�f݊����Τ j�.��g'ڛ�V{�޶�!��.
���u��	���B�#���]��>���/C���O_.pc�I�h�G������|�|=�T��Fĝ���V��.��"]���Y�f7�S�2,?>Yuf��E�	���>�����^1��Ǧmɓ���6�Z������ϕ�`��5����\�m�do0q�/���p����F�V�=�@�}�3J�-�ծ(0�\VZ��"�� %��xEWjv��zn�Y~�y�E�>i=ޫW��Rp�+TYwR:<��א�\?0�0�U!L��N�5$�\��a��j�G�uq�����B���F��3@
]d?% ,���²��Z�	��k�J�;�QM�.P���l4yn��wC�w� �(7-�`��(��&����?3v��a ���faf��z��|��p�׻��T5#a�b�`��)A�Y���U�0zP���/a�\y�å�R�^�íl�⅂.�#,e�3e��A�l�3o��3�;�v������ke!{ ��W�1�~�?UNX�d����V%�/N���ׄT��ϡP�g$�d],(�wn�������6�?Fm\�~\b�
���>/p��$��3k1QU�� ,����p=O�*>q��h�a+�#����7�Nn����T�;c]%ǹ��c���s8��= �'���x��i����V������Ђ�"��A�9tBCO>|>tƳY��n�9,�S�
[��"uaמQ�so��Z��ƫs5�~2_z~�����g�pQ��p�5E
���Ԥ
�	D����R�����h`�4��FJ`	ÿ��X��St@8�#01xz����<��Q� c���m6��IL�]�����ՠ��r4Є�~{���:��8���m^�R��0`����4�Ρ]B9�Y-,<�Y�O�
B �R>�J����p�|��|�2�Qx��@㮓2p�:d��F�F�*��|�������N�Sk(KX Gc|n'�n���ѵk���M����lJ��������S�8j$pa�"3yy7"�VUwZ��7�t�vw�H@4�v�7g'ޅ�|@�7�T�1�io	�x�:��F�0��´}doEJ�'p6\e������=vT�[tp�Ao ��ۗ�V��/��ݱ���4Փ ��TPI9|��;d��$%�)�G���Xi}j����0�?h�d���A�M�(����P�c�ůt�s]:Zƍ<Q�5V��Rh�����.�q*�'��@�Ձ暋e�*zG%3-�}O�dӝ`0,(��[@�2#J��IF6R��{�
ض@!P5����tJ��U�{?8:����Z��b/�i#��f���D�%�Γ[8*�!Yܫ� �
H�������b��p�/�/$N��3L�V��c� ��ܩ@t�OF�pS��K0� \����P��Ձp��̯Vh��|�3rZI�'ݒ1�t��'	S�І9��*,��/L��d��
��������[�c.�:�@�Dt���YI�����,������:���1�8�U���� b/'�t�c�g�-��ECY+��z�]p�\s� �x!��q�p�k�@>d5��3/N
�9���J�fc�&��Tix���׊I?w�G1~�Wn���,G�F%����nw��>������3
�"2��?`t����.���vɵ3�b��}���2�nZ�o2,��~r�z��#��]���jp�Db��W{�$��?���vI��:3��z<	pm%�\�{��M����
Eg_�pm�e���]cџ��]�*�Cr�jS {�~g�\\�O�zP:�(6~y�u��8��H���ͱ�(� .q��C2��E��|0�Ɲ-���,��U�N�!@�Na�a�R�h@�F�
w�b��ĈVc��p6K����6[��E��,��r���ق5�k�[0�yWc�a���L	�Rs���x�|�-AX9n䨚r9�� �g[7J�=_�c��=��UV����H����//���<?ҝL:9�;�U&�ɾ�blSK����$�o�tHo=��`2�}]4V�˶�.۫�8�]q����yA�0c9�o�},��٘	X�/q;s}����y�b�U+�3��B�@���վ
h?Ia�3�	�jcy��<�@����>p>E���XP�keM����%Eo�(��]��y�qM�A'j�:r���8��U����iS�ש�h<ڡȶb%Q�1�T�Mܵʕ8���+�8i�������~ӧOe��ti��7���i���	�cB=�Ŷ{A��)�7o&��KK]�b:ǈ=-��j�i
L)5� p+%��!r�b@O/��̈́<����t~Z�Q��y�V����
��@ѐ�Zl�,���&g�}��U�n���;c�W@�6Q{���*�ǩ,%�Y�s^�������P�z)��*�|")3�m`j��>�E��
����*2��c��(�I�߇y��a��S�S�Ƒ�龜�P����"M���g}̗�f�_���=6��|���L�,L򰳛�]�9zW�!e��)�>�'4F��]��_�Z��_8���Ed�:���Q`��������	W&�2+p"'7h.O�f�8��K�k�cz�F:=�8��cDD�ِ��5��>�i¤�y��I��P=􇲢�VX���fk�z��R��� ��*�U�0:�c�������r���K]��os����^���D�W��c��VB�G�l᭑>W~��rw������Te�Cu�������tŽ���<���u���iQ'`j�����=�u!5�\�n)���	
���l�.`eA)=��.z��Tp��^*L*Z&kMH$#��U��-Մ�3��R�l�g���)k�J@�,Z�o�#P�Q|�$��I�՛ӷ�z��������):h�*�/�X}�����i��O����6�zq��fq��^�W:�mQ�*0�p��o���v&�a����.Q
���_�����g49�6:PL���=A8@�p�֕�g�Y�,,d�K� l�Mi�����!,9��x��x�)I�J	m���*���#]�c6�YY(����7�Wv�復�~�d�I{�n�1;*ؙ�^�3�3�L�EUa�t�O�S���+^�9�#ǵ�c$�Jv�<�)1��?*��> �GE�����s�.l"�b4�?i�n���k��L� h]r�h�4���786tu���%��n8-W�QǦv�&�e��a����_�a�z���R	�s`��n�l����4�pEo� <��K�m/86�a��� v����NB�O�5^Ƭ$mx���Z򤏒"���Z���=����Հ�B�#{�>�߼���N���-��r�4�������ʹ�[a�����2@_pT��8}�&�i���K��7��?�g%�X*�b��h�u(uJZ���&��H?N��c/���=��F\Xb�5�5=tދt
nϷ^N������:s�プ�N��B{�R��9IZd��5"K��9�5.#o)���ݙ�������$zqq�m�$��{�FP��{��{^�y$�jI���+O���V],�`9[G����ť)�_�w��^u~�&��u
����%e�7�_� aB�8�	E���t�� Q�s��D*C����S?5�7��;�ڳ_5����c�:h��Y�Z�Ѓ������Ǭe�H��!P����=��)�\�8U�u��f�1Jk����c�m�4�W-\�z�ZH�۳��O!v=��*�.��&�9G6���g����B�`3��_���<�nTF��w��>nzkw���#� }/� �R��&��;#w���H��i���ە$�z)���d���QM�k@�����Lt%��P�|d���J�pr2�Ҟ-}��0I�E�5!�DH���� ��r��,��m���Jb]Z)�?B�h�-��Ö!)�(���>7��H"h��Уlw:M�ɤ�ВbSL�{^
��S�|�<��U
��`nR�๺��፩�-��!/Mׯ#+�E�h��+R&�Q���D���p���7m-av�i�����,�ϡ\r��8&�����p}D��桟T��g�J�ī������i���|2cD+�o�A����������ߋ\Qpp�L����X�J���!%6~�o�vK����.Kg[4�/ב1�_��ͥ�5Ii2�s�H���
6���jq.G�)�Y�d	�sgW�����e5��)��S'���0!��q���SN&FQ������Q*��G����!�@�x�Dy�}�)����k�]u�cp^�����u;a
�"��hn���o4C&7��֗P�[�4��A�S�妃���!C5�&Dc��?�/.+R8N`kjzd
�ѐfl�^<>�ل���u<��8q�ǯ�wER&�w��j��.�AE��<͇`,�x�՗���ݼ+k7[Y��4��.���?���k4����M�4/���p��6f7�K�::?IP#7��qn�63���Lp���ؔ{�b��`F�T5����P������#ڤR�9.� A�(+��_�IX��X�SOި��2;V��+X�JS]��PZӚ8�s���\��aE��h\`9��]r����-�+'�EK����cR���jM���9�Ae\�D�F�- �&MQ�7EVNw�ޜ��Cr��=Q|�_"FN�~!2��cl�Bѐ֊�:d���}�׸�C8^��Rڡ�v��L�D�	my�<�+�@�6+��^��`�f���RU��/Q�������d�'}�<��4\�d�@g��HH�����J�G�ҝ����%>��$1�o��V�F9?�>[��W��ا�_��a`Ʃ���d�VH��W���+��4�^K��`-t��qA��F�W�/2օ�`E�Q	;�
�N3�L1���|h��;¤�\�A��%�`:�y(fTF@�����s�`�?��:�Xm���P��;�Jz�Y�k�s�&�>��������bB�l2�32�aF�DIt��|:�D��)���jF��(�.�4��W�����	)V�w��T\˧�V��mOp�bZ	<�dA��V#��sC~߻�W����.q�"���:��}sd���<9.q��~%��(Hˑ0�o�$*��%)
)cک1T�9���h7��blivDe�U����=���U������s�ai,�X�B��ĎHYo�;���"]ڙ%�ΐr�ǁ�@�U5��p:���Q�7W4H�V~dc�9��~,~;���o؂�����Q���������2J�9X���%�[Gޠ�T1�ɗY�/1�����N�j�Ϡ�r�w���z/NZ5кo�)7Z&�!��I̼���X効/D���h���u����_�>#�%��iq4��ڴBO�y�ɻ3^i�,�s"0�r�"l��w�P&�H�A%4yMQӾhn@��3�_�}0��H����^�f�@ ��6*9�~�L/�c�9@��)jr_�,�K	�R��H�|��7)\
od�n�_H�#�\}u4�f�A~# H�X����%R�����m�"�S(��gL}�S1�!� n�z7�?/����ϟ�oP�a*4�1"��ń
�B*�*�3�����ĕ�}tfˆ��H6�g���xhų�~��s�)8|�H�%�Ănc���E����4�<"<��_�2e8��^�����?!VD������nM՗(&Q~H��d�n����
�:�cX��E�%�Y~�����~{e�3��}��lٰp�Q�3幥���)�k̐d������G��B���h�S�o5�S�Q�)b�pz�N�T%�l[�[�,��qmn���ɩ�ń
��*ӳ�jh�D����X� ���h�e������o\����K&SMX�}��ai��2��r�*kB6��v�����7$�>SI.	��^1F2譾)O����"���A�x���䣸��GTC 	�� p5csz2�pZ,�z�Pj*�w�����z&�NDPz�@%��Y�3H��0`D�[ �f/��F�Ϗ軕�a�K��l�͉@߬�!V\�u�r�뎁�N����\z�����: �^��B٥���M6b�%���w��f��r�N5X���@�9����������:Oٶ)���7sEp���iyWĳ�E����U��R�	�6�x���zMl���\������=����jK!`�騔ƈ�ŋd�Ó��޼��BZ� ^�yb|�C*��̴J�a4x��+	U�/�_����El��d��ւH�	zT�0t<�ud��W�l���X92RqR�$�YI�^R*/f�e`���G@��5!�dXm<N]�+�k̇J�\��E�W=!��ؗ��=�tq�P�xX�"f�~�_S�{�7v�J��S('|R=0�:����2=��Me�򩽜��A~��G�!��aBX{�{�˒�v�G���o`�����%��"��~u���)���(�H1!�Xo���/4-O��;lp��B��H@��/�{�G�h�ŠV&�vS��V�;Qf>Mݿ[�z�-������d�l,.^��g1x�}n��㕼קAYJ
^n��Ѹ	f���]Җ����w-u�?����V-kd�cQX�΂����2f��
EN���kB�L���E4%�ʃT{U�",^��Y�j�Ű*����>B�Û0U�������pĝ}�N~�{�{��aKK�Sl2�VS����h��Ԃ���kX�D���AR�@��]�V�nq�x�G����п��Ʈ8�l)�ƞ��ߍ'�'��V"�h��^p���Q�Q���r��A�?��H�T�\�[J�q�r�1W��,�w�1	�-vPE�e��Nwŭ^�Ö�s���,2���N�tH���FB��w�Lj��q�>$:�
]�r]f=���S7@�ޢ^����?�)��۫dz��0d���o��#��Ep��$ɫ�nǇ@�C�[��8�D�	s&�T�����}���I�*rk��&	/N#�mC����Y��VRq�t�{?sG���Q���_V���5'EZ�@����q=X@�е*�����Y��m��}�d��+~�f���(o�� ����M�,��;�0"��\0Ɔ�$�	yP��{F�gO�T��ޓ���que{��ɻ5O�8Ew@*�/��in�@o��=/�8�`����8�Zdv�tx9x���`�S�uI*�0�P#J1e�Z�]1gB�]��ä�z�-Fs��O�ɐP�n��E� ~�}���2��yy
�F�^(;�0��ETa��X����N����p�"�	�X�OC�.��]*-s�KBt�s���AļW~�D[-��Q	Yt��=�H�@ڑ��-R�TT�x�ɧ7-���z��sE<,8I�6�n2-5�)�"�gX|+Эiі��e�༭K�<�
�LCg�jT��͵��0�	<@�G<�_�t�͌/�Ν����=��J�I��J��e�5W�'T��v��m�ˍ�^�_�'f1Y��9Knvδ2~Љ��F����9�J��c���_�nĥ`��γ=�c	Q���7���g<o�R+S��
t#"�K�;e,����O�?[����'����x���ysy�-��T&ѷ7��_�$�F��7?�D	l\58��4�4�~v`�q��=�.g�����w�5������(�f�"�\Vh<Ya�2V]��#<ZC�P�H\��we��zhxJ9қ����$�i��p
��c@A��%�$�<O(���)���׮

���Gb����f6w�qS$j�q3[�����1I�<z�k�*���p�Ԓo��B�8�Į1��V��	�Ც���s�U�-V��e7�m�El���S��u)#q��QW�%��Haȼm�_��(�x��}��A����/<�*T|�/�� �� Ҟ���.�⥷��Q9kZ��I��u�ؒ�e� Xm*m������Ĉ' 2���|	�5�E$@��
{+#�c��q9�b(����T����N� ����݀�RGDn�]���k��lޭ�]8�(�Joxiौ��I�7>�@����Bɐ������AK;���2Lb�Vz�<�5}�:�宫���qݒ7<�j��I0��x�@��mlhF�o��d>��ĺn'e��m�7�#��}����}`��p�F�l��ϹEG�*zD�=�М�j�M����:�R)�k5A��.���L*��J�B�[]XEL�����e\b�ӏ�䞯S�ryX�Y�׏T��1�4��5�O���b����P���J�>ɮ���:ݒuT�͒�S����#b7d��W���xy��Cgr8�6�*��i�危�uyØ&�Wh}����u�����'Q�(<%4��~���Y�<:���b&|���C�/�Y��[�	YL��|`S����{8Yb`��6��Ƨ�z7$g���| �������O�v�cN��<;l��'�5�T0�(�4�c �EY��r�A�~MNw�π��r�{��m!h!%��~�t���[e�^b�"�hjs��X'~�Q`��r����~`W�1
r��2��I���-���j��ޱ�*�m;5[��_�%'.�$/�a�\`l����H�C���vϗ� �"$��Ǐ�M_Q�A�Q��l޷��-$��8��R�"�Ix�
�-��4��A��<lm�LQ�d�]�/넋X�̌_P�j�˄e4&Ӊ9�&���Ћ_~ٲf �*�t�n��Ee�3��y�C �&��������K)�+[v'�o�yj.��M�wl�Ȱ<�s�M���oa.A	Sq:l�x"����|�9�����ߋ{d�T>��MkY�/��NT��Y�7/ =�(tywR�:���u����D N�,�@��H�����FJOD�U1F�z��vRɡ�����%�9�-n@�tj�d�y9�E([�J���t0@K%m�g���\kv���`i�y�����FP��Ad��#��i@��298�z6��m���5�UϠ��k��P�<���$�7������/��?�TܨG�
@Dy�����ï�F[V�������D�7dim?�A�D�!+�9+������KB�� E�	��5+��cV�Xo�:'�ͦ����,���D��s�G _��<͜	��W.�����br�fp�m�����|�r�.���)��4�w���f����Y���\����0  |#W�>H33f��Y̬�Jl��Z@_�T�ŕ�-k�z�hv�",K�]ۇ�^'�abF7jGq���P���%zx�<�n��J6�󈍑F@3KT�^e�0�9"x�L��8��`�Ɍ�j���p��v��Lrl�-hL�?����,���e��5͏����?�}��}ʄ�0ӊ�4��5����/%����Oh"�� ^VH�!=����bI��*R7�[��������xc,����j�񲩳J�	�q2[�HR�M�%R-�A��9�[��w4�#~	 ���#Zs )��U����xn�Ã��e)�4��g3\/{��P�/%�|{��{�_N�=}����s����H��ҽ�5���-������jUQ�6��N�RoԖl^���1th�:!nG>�Ѭ��e|'��%uQNh\�ӕ�{ө��+aɃz_*� VZ�	�Ζx�ܫ1�v��I;ܯ1��+
��L� ���^�����?I4-),t�+nH����<h߈ayR�]ьRئ ��V��E��L=��v�Y��$�/�cA�G��.w��Zڴ/8�/�D����o�}AD��،L��~��	�N�����{�[��t�c�E?�u�-s3}%t�W� �(�2\��,5Iv3c�����?0�J�>S[�e:����*�l�gkB����$����3,�o#���E�Ҭ��h`�a��+��M*�Ƨ����&`!�r�k������)^�U���D�,J���2e<޶�z=b�5�<��/6�4NC��a�!���s�O��Q7�2��[�$���MyE���θ���ȯ9}�ι~��%C�B���� tO��H�/���|�����e��ԹP�i�Rgo4��_���x��~���!�\��ݐ���`��՚��H�ĝ�x#<�:M��bo������\<�[�_24�rY�����ړq��'Χ��_����Ņa�X��� �d�e���.v��1�IK�eUu�>;6�����
]�z���n)� F����r�-"B�+�k\�393��$~G��m���p<x��p��� ?(��H'�^�\��H�f���V; �"���p�J�+�-o���o*�'�r�S�D�Km�931&�< �v+�SD({K����c˨8�Idp�H衊����Xn�K��P~�lN	i��[7K��� �$���'�T.t��&uaO��-��<�,璍�?�%�:�5�R�I�?X�����cw��l�^���zZOM�����j�v �
��-�bV�ݚ y���2�'o�v�}��4���m����ۜBv{a
^��w���,�Lj�Q�����k�a��r�w$|��]!�(��0��1jA[�9�}�B�Wiz���iΦ~��-ػ�0 �+�o�$H��c�/B}���ի�в'hW��$)Wx��tj�"@���!��J"BNG�Ip�|P1e20_k�	� ��Ƣ�|�ׄ���L���A�}����+,y�^Hv��Dn����KMnKx����&#�(_�4�T�,���ΰ�U��nZ��w�G�G^�Y_?M����rM��=@r[?L��>%��+�S�����	D�6�,i�<�dj�&�>ZhQD�[���ד��8�9�;(@۬U�U�q��C�`���W������޳fb$U�N���m�@��o5�Ԕ�&�5f�W�M3p`$��Np�x	EE��Z���v�s���-6�ڪ�0w��5����r��vj "d+�M�v���}|��rg����u��x zb�T�D�LW�RN�pCbZC|����x���H�M9��YS�u$���Rp�-;A5v��	P �&�(3���V+�r8C����^���?:��4hR�w$���G��#D����±�!F;��F��&�r܅q�H�O��4G��mk}
�� ����*������Q�4��4���=Ĉ�K���z�D��"�5PH����K�{�6Vm�V+����
#VbD�½t�ފE�'R�֬k�fRĲK'�������U:�K-���*4	\��$�N���z�]��?omla��NA��BȜ7M˪n��}u`~YM}��W=�H����d{��~�q&[��RN�}@�e�.�xǍ��^�ZU<�uw7<����H�Y�.��:O,;B�At�|@��0u;��`3��Df
��Ш2����Iwh�B�m��B%� *�fAlZYWݱn�=�d�\�*�;5ql�g{��aȳ/p,7r�%Cs_���o��R.;�[ �!,3��xl���a_��F[��a�f$��ѓ:�ʋ�����ų_�%��W����T?��5� M�jw�ڙ�2��� e_��`�~���ݩ�.��Tλ^�qV��?:�"_��0��
�.�5��B�*#*�9pU�gg�@T���#�8�V��h!'��!O��q�S��6y�V.�k�D�	O?�X)m�۝��77�'(�S����J�����.X�R�Y�tz����D��h�k;�T>`Nȏ�!�+��PT�_Vi�]$�� x^���[���鐭,�9è�������?0�C'�x�v���\���Bɵ[�U�qI��l?T�Ζ�0K��(#˖!�crB/�!d%����:� �Ͷ�g~h͗��W�n�B�5;�ѽ͎{��.�,"9	un�#"e�/]N3ɊJg:I�����U`��$��k_$?��(7��Or��߶���ިs�^0U0P	PJ�J��)5��	_Sw����J�2�ux ]��s��+z�߃'�Ң�l�s8��Ttٕ'|Z�O���
�:�s^¶���?�ٵr���@i��*��'�B��3�v��T��RX�̳VY3�_r��:�@XR�L%��eM}X��Z��W��b{�C ����.�}�X¸=�DѨ`�R�n�ĝ�q�U�#Ѽ%ѝ�Zhi��Tj�AL.�|���-v=��jrn �7F僑��I
�[<��v�CR������ �|�}������ˮr�@S�h���ŅdR)�7C�f�W0lu:�]���e=�����F�rG=��e��.�Zͣ��S��3i�>��fwN_�k��ѿS�j���Y䥽ԨZc ����6�T�[��:��|�BԴY��D%�ǝ�9��Oq� ^b�f\�冬?�軓<�y���I��� �6��"�B*��2Ⱥ(j��Z�j6�5���� )��:;'�gǘ�?ԩ~Zh��Wʙ�����=�w���J��K���>�]��pAĨ�9���20H�xdt+c�F�\ ��ӡ�̰a�n�(�XG#&�	� ^ˢ���AHz;�M!���p�c�pa:���d`�N���a��U'e���ȅ�yG<Q���a圹p���s�s�6�*����/ޏ�;�D���TO���
~L&Uc��0*�c����r��	Ku�"l���/�`��QD
٣�����eD�T�!�FH9�A"�T���7�œ���$.6�� Z"ܡTqՋװ�h��3��)Ax>0,���dʧ�\%�j��?"_7*�eSQ��:�B�pɔ+c̛o_j�������w��,�K�LSȃh�D
�g����<K���%<A
�I#{����sL�M���뇳֏��J��a�P~��*.<S�9wx�x�Q�<��k�*	��9�ݏ�%).�WsG]�Nz^�`��@�>U��`'��\�d!���L��e�]+b{��y�dZbp��K�?����Yk�q.���II�1�y���&uG��y�N
����;S�Eߘy���۞^�78��E��d��b�槢�c�/����pf�/�
���q ȹ���\����ϙ�(H�R�'�xL�G[U�A�+�hN�L�e(���Kd�$k���J�?��J.�5����ڡBJR]�&�7�6Ć����G#z��C�ϐ
�%�*�h����S���d3�+&���'��-JU{	���)}�F��y���p���_5��e���U�'+u�%(�"%;��p����Xq����=�1ũ[��I�27_��+p=��(�6 ����ֿ�^����aq�F.<vh��U/�1@f���z���|{~Ed� �T�AT0�z(�6e�G�(�{m+����mcc��(�a��O��~N�d��}��L��ʘ�{�w��&'�'�	���9c��l�D�1g+�p~�%%��`0�`*Gc�T��R��e�`E5ꙶS/��5 ۋ�&����Պ��s��|���PE��k�� z�x����ҧ�_~�q�*��pk?�o:鹴��(-��X���tV�F=,A48���jds�@��E���F����&�{x¬���1�%�MJ �t��WJ��u�(0S�b��A[<68ĥ�� /=|}Ҭ5���~>�q�"��BJ�7��#��vZ�oMԽ{(�QKДӜ,_�K˷����]W"I�K��cpU����C�E@=����CJ�|<��\绲J�!O
���K��o��|�]�D��	EG��a<�Z���8� �nu�X 9t�{j�(�����F����8K# �`�����sv\[>�z�.���.��-Jĩ+��J�^f�١�]{��+�R�Í6����'$��|jv�����Y�x�C��t�������ꃓ��U�^��f��<��t\pj���}[N����V]����|��;�p� ́���I� �=>��!AS�.���)h���Ya��Δ��F��O'1 a���Ʋ髻ZNtGғ�%熒F|J��8��@�\��O�����E��Hx�0��1�M�D�~�51�ϼ3�6A��PN
Y�*� �E��B�v� �u�����N��-�q��ځ�!\��i Y��x���`�вf0����0>ǌ��]uSU���r�䍾9#��z�-V�\Qӄ@��i�Dn���~�u;�ŏT��l����GT�h6U����e2	}|+���$?�M�r��A���휂�2�%*�����n��T�q;��$���e�j��@�r����*~���������XC���S��+ۅ�Zl�WM<�(�Q6�j��XQ��Ԓ�b�/V!P��:U�*�r�c㜹Ä��@��"����R
^&���gK*A܌�{�����Y��P���%��ܶ,��]#�bR�NK����F�8k9M�ܟn�
v��-h!?�s�W0�X>0π9\�(�����y-
%Hu�9�z,��D!�~�w������s�Z�b6�-Q�Y^Fa#���}qj��FV�;���rv #��@yH0.�T�Uӳԧ�I��T��~�见i2	:�g��ܘ�����5R(J]I���$���Z"��+d��>��Za'pk��Q]�)����Ceg�;� �N\�#X��+3����H�X�U$��a���i�$�ۈ3��%>Gls�o�N�-�U�G�{��U)1pˣ�H��:'O$-{��5��s/]�)?%!6�g����þv��B����CQ��t��g���h�/�X�]�3MT�T��ss4'p�^��rc����7��R<?���v�k�.H�}n���|8Kï�B�s>����E7�Q�&�k�\%�2V���>�h�@�s{.���k�~�t�\@��Sڟ¥δ�I�ˤy�T;�&� 7��l�����\	r+�}��h�f!S��P�m)g�b���<�䚍(?B��Q�}8Vs���zU&�gcl*����Eh8mfG�q+/Ν�0B�>L��Lg$>I�q����4a1�c�~�]H�j��y���B/��w�,��-��[�y͉�V�T��՘¢�K).,�Mq��X��%+���ጺlآq���B~��|BZu���<���p��f6�f�p���B�5��@�$��	Wo^��ȷbB}�f4�.˾LXEq-,�iZ�M����c�y�|}s�^�JALbW<3���t�m��3�ω)�CQ��W��k�}��T�w��#AZ��i?4yz�w:!c~��&�Bh�����Ϸ�d�6�|L��<a�~��v7���0%S+:t���:+RK�`zV�^����Iu��C����c�_���±����Q���G�C
��)��������k{%n��uAն�2t��/v\�4���^uf��c޹L;��������ŸL8�����Y����\=�>'a�'59P
(�-�����NX��������-^N�ɭxv�����!�s�^!���:d��*�f��Ln%�2@��	���^V��W��g?�/r8�/�G>e�R̎�Qt5k��2��y�+�J��ҳ4��9 �0��K(	�Լ:�i9bi�����K���DEt�!C?.�G=��S����
�n�V��*4<B�E�Һ,H��,�����[r���$��f7�HN�/����e�ƭK�/���f�LM�����M��`i0�$F;�n��c����d�,_~ ����ώ+���������~8�g��$�b�g�f��E�ւK:��B����O�6�#�Z�I�t(�0��9hJ��`�X�/�XR#<�t�R��l#=��	���ɡ�EMH�z5��
]��{ve.�ƊpS����si9����*�@I<:��Ͻ�T,��Z��(�U��ꩃ��$��qq�\Q��T��]�O�C�$v�iꆜ� �k�����yY���t1���h�A�L+���mb�;��B,�-f�&q^[h~~�l��%�M��]�cYR����͸'fz-˵����ב�6+ew�����]3㋜�(x{��8F���=5�Q�e2u��;Cִx����WW�)�|G�=���0c��S9�lς�Ə�P�1�u&��Bi�S�C�ҹp��Β�aCc2F�t���:���d&=���( Iv2N�zfHcg�_��Wɝ��F\oO��m%�u(YWL|u�)���)�7�y/ [��*�2��"��[��H�g& �N�H|
wL�Jg����<=�L������3N�虻�ǋK�J�?���z�&-�<C�b8��V���d6r.}�������[(������I�&��۷�����_̵��V�.y+��	r1�&�����ꌸ��Qb�t�I=X�*����yxX<�"}��A��ٱ枾�Gm<s�x�9�Zq��8F4c$= �6�e����қ�y��ɇ���E�8�k��e�m5�f�2��x�{P'��қN��	�&��F��,~+}阶�8-�҆��Y}��`?�=7n���Ҍ��GHz$n���l�,0Q
��Zx^��;�T�
��,Uv7X��w��C��Nx��l�Q�֩@�Ff�R��h��	�J ~�7D�=P�\���.XJre�P��!$h��P�=����U9.Ɍ't�KN�Gf�@�����!��F<U3 ��f},��d��Z�B���:�ۦ�0:S��-������(r �b�(�O��3��d�Ft�iW�J�-؅͗U�t;>|xN�S�A*����K�#L�Q�vU��j���i^�@�Z-!h��kl�73F�D�u����t�etKಪ��8�˹�	i�X��^���\*�'ܫ���M�9�rͨ&ẖ�=�<�d����	]ܪ�随?��<i�P>�L L��hm��ɉ��j���_ �#g�~��)�s�{j�Юިd���!� �[�r�x8�T?� �8��bF]/�>5�bB�A���GO:�n@���"8�p�E���8/�\
����2@R���Dg� �0�K!�x&��]vE��q��v�e[,���Nec��Yg� ����7qA����Λ�q����J�����*+�&`��u�>8r��NTF],��N(�g����s2��������d$Z9`
R��۞��ƪ�+��Sg��ݎ�@#y�I�#��U�5��Q���;"Q�����T��c�S��o�%��/d�溚M�U�� �Կ�u'±�v���/�cE�*@%�7�+�rf��\�ޙ�h_s�F[�&K�3.�&�b�Є��p��K��h�,�0����a�[�ݜ[���Z�{���n|R�di�N�K0_6��~�D�s<X�awB5��1��P��+�(�����l���6`B�S��®�!wd����>M˛�`���^#�)��t#��r�k�ٲ��|��f�Q׏�$EƂ8��."Lv]����l5�˜%�d�
��朼� ]�3��k,�3�S��cI�^U�B��N�G��1��>顓��%z�����7���bq���,�E�G_�HPM��RN&�Ȏ`�����q����*'�����#ɒ�0&��9�2HB��T�f{�k%2~Soj�<?����k����2�2��o��"-�w�������{!��0���g�	Y�myq1�[Q�U>����%��j��B��]�$�!$z�@|x�zu{PE_`:;�12h�X�������X�d�s����Ҹ��7�8�6��ǀ4:�k6$�s'�k$q������C��UC
nP�[]�J����)9�Oȑ�>C��A�P�����5�#)����vMl���9�,���D�[�|�oY��Ln�*��ڕ���T+&r���
5q�x���/�j�!Sm��徭�'�BO�l����j�-@��i��.]U��/��hHxd��= �л\e��� ��5� ��b�r�qq��a����UCI'm����֕M-�(U֙!�KrDh��K��kf�bm^=/�3e�?�˴*�&ȣ	"cJqq�:_�>��.��)�����%�(�Q�%������qOC�'��ʞ�*��o�+7����Q5CY�/G\"h�z$L���5�,��߇���C~�3��V[�P�U�P�y�������I4��~��@?9]���&EU�y��=�(�Jm�*����n~�W倲J+��Ʉ�@k=���Ŭ�7yG��']A������8����L�r0K��4�¨���|e19�&+m�0�J��i:��ɠjJ×�^җ��S[صv
�S�Ӵ8�Hw�g*��Z&���b�?7WE�[�<!���2xW�q�K�^
S���h<��x����Ę�\�wb�֣ �D��Q�݃e�����}�	��M]Ȕ���e"�)�-a�3s�(���s���ns��/�p��Uc���&lu���%�-�ť�g�h?>��&�?)a�m�{	��6�{r9��q�l%����f4G�z��<#�Bꯝb�Jj�����0���	�	-���z9d��j�ʱ�è~���W�D�G�]j�F���p�53�dZ����8=��3X��s6-Ɉ?����5�O�<s��M*��å�H�4�ߢIY������̳�o'"��T��<�"���Q=,$l�()H�MJl�(�����<��Q5�8R�4�+ZC��#DEz����iV=�~c�ri��}4��Й���s�A��iB����z)�2�������!��HZ����D��y�<`�X7�D��j�kE��b qަ"_�\�lYm5�+y�>Fk��-z℠E
�|"�+�y�+�!n(	V�� ��Q�Nj���[�S�p�Ɏnj"�؎��S�c����)JʙT:�)��|���������(f#�2�N���Yj�b��U/k��\u'E:�K�V�>�Jd����K�B<7],j��r��1N�_+h�i�5� ~��A��{�D���&�'t|G���@Iip9+eFy���r�C�qv�M���Uzo����%�i��8���e�E 7�s�1<�NY큀�r��ۻ�w��݀W���[s�g$pz�j�m�f)q�s:^%�4Λ��[��z댤��=R��b�R4ϪRAX��[K�ZM-�]�A�����C2�'��A9�'H5�u�H#k������3�����|�矄Ȧ��#��eA�5Xf��Y,��Jҗ�
݄� �r1��wH�!��w����	� ��<b'������l�C�sa��e��-V�,��|�5x����gc�D@eւ�0Z��&:����d*��[�c�H�i:\TǺ���$�� �_:�	�R��H�s���d��2�Mב-��@��4i�!�vm����þ���<7( {n'h�Y��X���G�O*����ķ���l��}�Rq�.�tc͒��䁞��`�+�������1/bv� �ʣ6]�N�]_�o1(�_s�/��|-��,��DDp�U�b͋v����	 �o��=����kh��#����d�:Gꖦ�A%D+��y��"��Q��
��T���;W��ҀǦV��qg�mٴ�����UH�%��� ����F���n����jo��d��g8�|wf=9�����]��؇'��6�=
6[F������P�[I�魿�J3v#�ؒ������#%�_�B;gSS[F���)֋�3z+5��/l?C����'�l���O��Y~w��D�D��f�N���������f	ʈ�ӂ!���y�m2:]_+�f���ৈA[�X�n�p��֒�������t�o�{�A�~���Xx�o/�TB!�E�L�����C���~�:�￪���Y�p،�һ
-(Sf�m�逭���6�������|��9?+�@]���y*E�}_��ο�.=(_4?S7J�淌j~��ʃo��"U1K�_�ӏ��<)���䠥�\ֽۈߓ���iu@��{���,$�d1~{�J+EcĢ;;+L�]О;��1�0xL�Gh�wD�l<�f{3j_#H�@�1-�;���;������񀠄��3�܁&_�m�X.�֋Ae@��2*:>0�SB��}#JK�w� �&J�i���n֪�$����o��Y�ۺ7w�_���`:��f���OI�Q<�$�C��3�^V�(�/I��ye{��<�j��ǫ�ڌA��0�1t��q� �=�5G{AL��((���+�q��>�=�d@W.s��PH��k#FU�b�п��A��,P�9n�����5�eY,�%�VM�&a�~{U�o�d��+$/�"�����kxt^z�v����޲�3TR�iI��f���������4]��=~\H���^�Z/��x~��Ԏ�&�Th���hܯ{���I�k�z%����x���z(XGH��H�U��mW
��b&c�A�G)�a�D~F�n\{mb��,��&�9�Dj��eՏ =/mSI������͠���F�jM$�*R�e�Js9H�l�>"�&ם#ds.�D�L��e��Oٖȫ�l���G���S��8� �'N��Ҕ��8�9�{�&2U" W�6�|�;)�"��³ƫbN�#�&H�ʉw�٬�؂���Y~?��!,�A��!18l���DG�.e���E24�f@e�$p�z� -/��ztDY%�4����_�t&/t8�}wƤ"��4��8�3��[y�3���}A@Զ#1�mI��?�̣�����,��@��X����Pm[JW�����w��f��7;��g�?�҇z����dI�H�Hg��r��F�O��*E�\��S+�\�peB��\�..�7FJ���������u폢'��o���]�����U[���Eڀ���٪�&���8,�db���FB�DЧ�i�߽�u쉶h�����g�/NxM����;��~�6��gM�<w��D^�.����<�u	����92�E�k���k�O�l����<��r��t��<�U���3��]pD�W�� Q�B1�fѩt
���&RBjK[�1*��:eǔ�@5�.)��9LU	E���pl�8�}�0�`��ޑ��%#_?��a{xO�\p�L����ɓ泌@���r��l���:Ĝv8��.���c3�չ���0�cR�U)2�B��3OفZ�j%)�?����h����M]{�����SX{Ǯ�~��m���i�H5*_�r��W���l��D'}L��nϘ�t���`������[�m-�7ׄY撞�z8�C#2چ���-�$?W�x�|�O�n]�ߊ�G��6W�"U��o�vh!$���������s�tIb�� �Q3�}��:�}gc����e�M����W�Ѭ5b)���&��*��Mwp+�}����ޢ���:�]�j#�&QLJ�\�[�C�`p$�W���ӝ�e���X�Ɲd�$ �_�ݨ��l_v5�����`��7�^ͧ7O�i� RI���~k���"c���Ɣ���	��ʪf���Sh[�#����z��/�yMD��kd:��j�����uJ����C�H��I��~�A]���Ab��SD/�m�<�\O�#�d�8kD�'�{���Q��S �j����Пy��?�����	���
�khV<ABs��*�d��My�5u��W�6,L��4F������U�ov[&��h"tD���1>xe�����K�PQ�c�4w0��x��Z���f����K�E ��ظ�N,,5�����,*ƾ7����!Z}�7*Ci	hߐ~(܋ ٲ�^�#���?�r#�2���#Oh��%�ar���������r���q��u�:��{�,���X~��׳L����j�7y�"�q���0���튅~��E�M�s �j��)!�zw���6����ڪ{B��\���r��W�s�m��˦�������O;k�>e��crD8��{(��XpH�Q��ZX+۪o9ҋ{�q�[K���@-�s��vW�`uI;���y5}�O�;0��6���������@�v��]"Ж��#없��(��It�Y>��[��p<��E��G4ZgR�
�^N�o5�}p��;?�6��������L�]>E�qд�9�2oMGOR[�.:��m�á�0-\��y�m�K4s�V� � f��D��S"���eC�n;��q�����.�f[ЭD��Z$w���N֋�lh�h$m��i���ӡ7S>cP(s+s�[��9��T�[f,�������"�ϛ�q�����K̏@���Qc-q�- bt��Xm��ޙ��{&3�����d��u7���/W���k���o]���#�
���t:@���Y0y"u��O ��w��R��V=��1|�ӃY�B�%������±+�z��3W:�_�轮;�Z2_�*#X�]��������8=�>��;�\��D����OiU#���%�; Ξ������R֢��<Y���9u��W�P
�Yk{�o�@����@�j.^�����9�����~m�O��5�9�+��/#����g�)��C�jU\�;R�ҤG
�Ǝ�_�qP{,l�R�EH���w�w�
��wMA,��2�eZk�P2:��ة��ޗK�w�Ñ�I|m�h�1�rw3b�Ҍr?[Tф�:������[�}�G�?1� l��`
���*=��r48��%ߋ�9�%�=�������|��ߑ���X5=��M' �C����M�j�w��8t�Vu�gY�-
y�7�6z�PF	�qw��P4�[�-����'o�����})��y��8C��T�qX] �D��:$�В�b�?���KBQ����$�u�OD�ق%�p@�F�@b��6,c�:v �F0A�y'iR.^��-�l���y�' Ji���;�Ust��s4<� 5#j�2����=����݈!�'�m�`�Kbr Ѐ'��X�&�����B�BR��=���~l<@<^��Mm�a���$��p>~D���.����]8�a�M��}�9�tf�Bh�vPа��@�:��͉��V(�7kTo���OT9/�ʥ��G�
����"�Ȥ��M�o�b��N�8L�1��z?�D���#�x���ӞR%	���I��ɶ��|���A���(�n�FL8�b�Ύ=e�/�Ө�02a����FR�t;Ԟ�K{��I�������� ˖�����D�������/m�Q̋��iJSc�?]/�h����V��֘H�w(��fvUosA��P~;�{���-�2�����N����1�᭫�p4���Q����o����<� �-�h�3c�@w��_n�¦�3||���mr�����_����'V�%B@0 d��U)���c�1N��p�i�y����}2�d70���%J�٦8R���[5��+�a�rZ���!�f1#;��>H/�[v4?"݊Ea��փw�<%M���v�]'�ԙ��Q��g���-����� S�d�-=�_��Hv5d9���0�a�zUz<(_W���Q�)�+�m�����y'h�z�>A�''H]3�`�3�A��l�����U���8��H�hM?yX�ͤ�1�]ۓ,�$��VK&,���a����w�~��7�����}:����Ż���n�}�3�z�˺z��H���eF��E�[�\}����ܤ�B������!h��~6�y̤̖Wf^fȚ�`L��lv�QW�y����C���+d�I�P�n����]-#<�Eh�1b�E{�Y�n�'��W��e.r2`,<,�p`���S�2*��������L��z7� �b�&��B�uK�ɱX6��d�5�*�M4�u�]�7��#�p��%م��f�!:�Ͻ�+-�"�H�����&���)I���-���#+��sx�y�����@��7�+�ں뼕	�����Y����F���v�N��S<P���-�tx�	}�5��M#ê�#�s����+���sj���H�<C2�Z�i�؛;���}R��	�ao�G��.oO������M�������-Ѣ�돤�6iYvu�"m|ecON�rK�s��2G
�V�`w�Ҭ�J"�3أ �x�I;p_'c�)��J=UL�o^�"MNT��M�d�Ch�C_�LB��/U;��a����v�▹�g�~R�a���-���U�̦��2S�ѡǴM���%����!p�m��M��Q"�V�uM��9�	#�GRx���S^c����m�������R�k�"Χ~���Kb��f���WD5R
<��\�%|;e"g�ȼ�Nt���۶��cs�<"!�H�Hiec"�&�s�b2��7���A1R��8A���:	�8G�����i�9�Ԫ�V�eB��!��C�YO�P�@%Q�vN���x!�e�!��V(ɧcX��P�K��#M=�(��j2�g&�@zq��6yQ�z:J��)��3W�_�h�^�ze��\? *#�uD,��[����D���t��k��2�8���q�H��s�f��V`-����/�����K��$�9Q�]��v��J�(HVxjc�	��f}b�5e����}�����А�K,�$�E+���~8Bx����Fl�sc  M�t�h[1s	���{�C>/��M���W�.��q0~nC30�M�M��qb󎃘���zT*+dcHD/�UQ&(�2�<���+��	����KO3-i����9`�3F�~��a��O�L���I�g'�D�uñ�����]C��̂��;���#:�i�Z�ߚ��L�TΤ��mPďeD�ٌ��>��M"�w�k��F�?b_�wT��Gέ�
��3!ė;s�I�û�:'�KV/��n��������Ơ_��p��w��Pc�/�;�DQ��\��q�5h؜�C��B��{Z�Q�
{����t��g�8��- �g;�e��s�iӅ\�N��CX;`;�vY��9���wu0��-\�$7\�?b\���Di���K}|,}aP���7�p�_|m��8J��g�0���54���y ��I�f
�D_�Z��h�:(�m%�޵��d;��I�N#��{Ԥ?#�j���7U����lK�H i*��]>�R��\N�;�e��WF��m�{���I=xh�)�3���V�tkM�+���ՠ\�3"yD�����@dV\A+I�;�_�����L���b]9USZ9�D�ݡ�ckg\�z�[�٘�vGuRL��o��ζ3.CG�X�����i���䷶�GN*"X-8.C7{�!a���x:+Z��O�S�9�kX�x� `B͎'�M����L�Ӛ,v� 2nA&[ �ӍE�hZ�W��M�=��I�H8l��_����,�5椬b�z�#8�k�M��j���j#�w��͓��H��1#�8+y�P�T;] p/_Ɍ��OU�_���pQ��8}���qؙ33G_^@�~x�IZ��m���߆H�������S�%��˳����Z��|��v���=���?K���*��Ug4`R�]Er>@�c��B4L������M��o��2O�꣎�H��.[�(3zl��5�ԁ�W����+X��"�I9Ԋ+�]<\Q���C�sCd��u��X}����w��w"wuv<���k����%T���=#Y�	.k�N���+G�)�|��#�{�e�mW��EIv�:�TF�,	+o4��"v��z+Wyv�	���u����@�%ee��F/y�C���A�t6\�R�G��#��Ru�į�N�����t�ʫ�ot�YF����}�� ��,�@�����tDc�"�˖x6�r�{`6Wr�R�/R#d�GnQ�\� �:�1���Y�q+ƫ�C�1*�ۜՌWvu`N�&��{]Z}�z�1ɪ4Ʒ<�mB�tl����9��'��^ߩ��j�:
mH��r�5z�j*Upߧ�ʍ��Q��-u8'��wC*���iX�x/���`���υM�����ȕ-$�4 ��uI#zc9��?�^k�#'�k� p:h�+*�p��Q�(�~�B�:>Ͻ�g�n�b�QO(��+���8٠�G	�G��{�*�����A�ȷ3+����#5z�Ҹ��6�b0��(�2Ivh!N[nV~�9!��h���᯸�����Z�$/�I-1@_[����p#L���$��jK=ӫɷ�>��./n�ؙs�����=ؙl,��/� ̝���J��#r^|����{yQ�8qj[��S�P4X��Ht9G�3h���㕒�e�T,.��-o���G�Հ�k�ܗA��5�����ʌ��_���Pm�`�Z��P��;��M��Ej�$]�@234nE��M���0_���=��W��4�p�|��,.b���(�$�:cC|�����w����0D�G�j�0f�7�Ĉ]��8�4���h����n>�3'�0��]����7`(�
��0Yh&�>SPT����T��͓XЌf]Z������@����ވ��:�qf%�X<yÏ�KO5,�D��L�)D��(�H�����G��{q��&�IJ�	S��9C��%J�WNQ��H\U,�I$���{%=^+���������B/�K�f91T����8$�]+�i�w�����K�ݢC�t�u;��Y�k���T0W�/���a�h7fW7��Da��]�ƈ����R^-ߨ�K�D��ۣ�ڲ��ҭ=i$u�N'�Z�<�%zL������y���A.��3>
��kѴ�jH�Uv�vE�r2�O���e~����KQNrя�,������hJ����#�����Yg��m�bD��c5�b���P�L��#�'E؈�M�`����1�Ǩ+����Pfo��_�ց-.��	���y���oPí̊N�	�6�R���Tb�?c>ڽ\��(}ᨠme��S�D�C~�]�\s���`�iA�Bqx��Y}4X�Fק��� ��/�˓���~�����V��U.m�
]�xl�H�
u��E���B�"m�"������]��k�.;<-e
�*�O�Zl�� ��ps=Ī�g����k��֔V��y��"0�����
�}*j9��L�'��a�yf>����L,r��cʝOm7#Q?��W�W��"�?�4��US�OE3d+(b�dnT	Ax>o��,7�5^<�r 	�Z��C_peC>�c��?y�}�n�����0�����>�P��m1s�ݙ��ٞ�˩�j� ��8t�Y�<�/E�h�A��%�$_��E�c�ҪJ�����X�Lb�}��k�;��ݶCaVLH_�
����m�°��IC&�8�P]�X�J�o�D�=�!7�.>3�x1�i3DZ+���T���_��9K��M��}�?�DI����2HQ\R"�� ������s��$L��ڐ��"#�U�z�ҽ�y=�4{Gڼ��(�9��;�R���vv]���bp6�u8Q�#��>�L�y\�~ɠ�=P$�դ��i�˅H����,\G��k��@��Z�x[X�c baP�l|�$ER`˭~������a*�c����FZ��v�����n�9б283d�
/�:&-x��nh���%���~�y~c�<���Dh��R:;Zr�4Rt���@<&bk��D���8%?�}�G�\�!>x���s��1�f%?��)�	�f�fH�ɳN`�e/�m3
"݃{����6�h~*���v��Z�*����U���Bv��;`6b�īlC�:^ig�M�oD�eV
q��M]אV��:�a����~?�E	"���z�v%Bӌ��q��[����t��eyy��@Q�Q�~Qs�L����*{	����tӣhO�Ϥ+�D�����T�\'�7a�����^uG���H�܅z�V����0}�a$��c��r��^j��sX�r���)���[�;J`k\t���� ��h"���RY�3XD����:�ϳ;�a$��ˀ���:�]F?�'�X����y�����J��`���"{l^���mz���"�`=U�S'�"�S+��l�{D�v�7mV�^AT��7d7H`6Rw�S�����-l�>hPЍ��Ę썠d�=˽�c��Τ�5F�d����M]��R>lң�#@]�����{^�r���iR��oMըN%���O*���wP>Y�&f'3U!_�n�����$��mwz�c�X�G�Q�u���`ya��ܺ�ִ@���1R��,&�:��!a����1��x@7�� z�]Sg����GI��ֆfy�*R�*�=@�a�4l*���*=��:�(].>hJ:�M6��*m�7	:�"dGx���zh*' `�r�����*�´t8�Ǒ�jO��$�2���+���)���:8�%�; ��"����K �ke��d��<5sI洉=�-[#ގ��t{m��D��83�"%�ղM��9F�R'�؉��&�N�n�$iG��U+kyn������QխV��<���O�0���͂ā�=q���yF;d~.��Jjͱ�z3���. ��!d�� ħ���n��o�/��`N?�������v�S���O��~���0������Q���6#J��W��5<:)'S�q���I��R��K
�Fs���[�j9���#����m�H�^;�mtBi�uX; 	m(��d�@�J���lAޓ]�t_��.С$0#�8��)j��2�B�+_S� _����GM�R����	��n��l���u��Ǒ"�!�1�ڟ���L� �5�~t��G]mL��O.��$�!iL�_u_��	M�'S��9E��,�B9n:�`y����~�m$�)��/�?��p�T�r�r�3p��?�����C����KI0��N͒�g��6�� Ҵ/r��I&j�8�<�QQ�ЋJ>]{����4�5���S��,�AA���u=�����-C6v�b��_����S���/����e�\v����-�
�e����2oob�8>4V{�&��54�=�Y��ܬK���L��P-��q�K�<ܷ&h0�����񣖲���{+��<�`��A�A�
˵8�m��
�1����%�~̩��&�J�}�sϊ���.ϳv�6�ݨ6��fR�'[���{�T
l��oOY���<��r����fr�ڏ�M����O�4�5�W������S��M�T
�����\1�z��?2�tK3�4�˱�����ay!S�{U+tN�r�o�+�[�.�f˛�7T[I�$ԉ!�2��8_yF�]Ȗ��nU6;�u�V��Ȝ�Hm$��Wj�t�.�0���jr�Ddc�wt;�(n�d�4�Ԗ�^�Ȣ��=
oެGw��uP�-�{5�0��<�ƒ����z93�Wt�8"��䜫#f���v��qh���M��:V� hw����Wі�1b�њ�5�,6�Ǳ��Y)��EQ�_7��D���0�\�a��d�&u�éxn��;��*�׾�b2��A�*&�G�[C�7���2�W��I�~��\�Y{���xD�UB�`R�����&%	e�|�*^k���D����I=0O!b"`�|T <^�PZ��U�Zx�ɓM�i�Ы��7�tfb{�w
x� ~��f���~F��W1),��5잤�*2�>��t���x�2�(��:���ޢ�u#N�l�K�j�V���J
5�>�fM)x���(z��$��Z����r��1F��[��O'R_Ƈ�3 9v�#�;��5�������Q�lT��e'�r���=�#l'�mc�6Jm\�F�},��
��������j�U!��ں�^�qS�a'j�0I�Ȩ�Hɨ{��3�H������ߍMz��������t��.wA��c`��8�B�|�j��f�Xi�;���mU�����L�.�:�*�ܡ�2*��h#�-�O">vE`��	�*=��X!����Yl�:;�6Я;�E���(:�{,�/�_�	��k�q�ٹ# �9%6�;���W��i$]���&�-X��k��d��Z'|�aWڹ��Z��>\.�޸^��g��A�����'w7��a6[c�V��C��G.�x��H�y�-ei��lq|p�kFث����YH������e�u���[]EWZ�1�5��Ll����Hs��s��u���+C��x\*.-�����N��'\g���4D���fU���!�.F�J��[�$��H�׽����^R��!�۬��C������E�i7��>ﬦ�}�ܬ�:h�"J�^r���#��QZ�q��ھ1!?+����&9v)5&KҞ��)>���:�0���Y!��(1������{>���k�-�c7*������>���_cSQ��?=T�T7:^�5��\w��Gֆ"�w�j��1]�����(?!�C}(j���Rˊ��|���=v�LȲEj�&}C����m�ϯ�<�X,�4*'>�?]���̃��Jf�#H2i`!\��7?���	�V�N�
��������׷���B��jE��s[��ﾜ)�G�tS�؟����w��xUIӲ{��[�IT��ˡ���|l��x���ܿ�PE�[Z�J���{�)Ԗ�bD��;q`���*<�ɉ�$������x���$�Mf�����|X��p�^@0"Y�ǒ�bJ��e3����j��������]�p�w+��8a5����-:U�I��w�g��B.I�ˣP����	nڇ��U_jA��G�ޗt�(6?��N�r�y����h�X�
3��"oS���A�n�	���YWu�9�FM R7w�9鎠�|2��uy.�.�ZP��"Y��J`��Q�[7E����;z}܉�j+���.�v�kE�.��cj�3>;|�ɤ�i��Q@�N���"���'�q��~1[������B0zF��M�_J�:��{�s y��&�쾟�	EĚ9u�o���ś۸�K:2�����sn!ca4�r�S~�U�؟�ɺ�"?
$޸�`?����"F@��޷9�ɏ��γD&{�]b\����`�e�\�Pb������RG��i׸�>�h��vE�J�/���]�V�{�'\��c<ӷ�nH��e�Q��߸�N	��_PpY��v��a�d�<`��0��N�<�g7��i�6���oS��y�_�v�{��ùz7�Ｊ��Kn�n�
�y_H��yƘ7�Z��Cb인4$��%)s֒���?}�;�	�1ٳ���a4��̨�8�P �4�aӐ���X��V"׌�g���8��� +A�r�6ʮJG��!����"���-�[Q���H��e�3�ί��Y��Τ���t��k�S�V�+$�Y�/ý�K[kL4��@|Z�q�WZ�XZ4�枳�
U��sFd��/�:Xgz����l��
G7��p�ͪ�Jz�y��c)):NpqX�
�2�qX���\�� ��6���� ���y?�{�+O0���L��u���h��_(�/���Ѯ�m���ߘ�	��.��q�|�?���S�nO.��&}��C�>�մ�����/̻�㺐H��&��zG�u�k��H-�]�-n׾�v��xF��e_}[쁝����!P�"��.R�J�?�b�[��7L��5\���$�t�D�xV`�ۤ�b4ѫ���G	6="���Л9����ȶ�Y%������pM��i#�[� ���Z"��:V&��f7"p~U�g�yY2}N�37�u�W�.j�j�:�u�:Az���]v{sLb��L��:�T��?#�q�T})mɸ��"�K���� O���d����%>ߤ}���*ŗͦ����1ڜ�����%R��J�����7�,	'���g%��6J��b����q�'��TʒV��ݛ4���*t�oM�0�_2!��>��8'3Ng� 
ro��QD��K�6~�1����:J�!,_�w�:�|���M���~���'��N
Tnf��K��,P����r4�|Sݞ���oQ���lr��c����V�bJCD.Z� ->\�0bW/%Iͷр~/�o챍b}��:���/A��9�@	�"��O'�!�j��N{#��UoG�v�?�{)�E���Aj�a��OV,n�2t0���|���I
M*��k���b`�a¥�k*&᠕S-���~<gI����f%Q�_�~��X����a�C����|A'�p����K���=��Nɽ ,�e �����O�Q�"�2�	{�q�{S���giI�C�e�C���j�=���d�v�;䆜�)��Р��
��%멕н�8���3��1ד=�Y���_�۴�G�8a��N�9�O�V�nٷ\Y�O�{�5^5�s��M���� ����N,�͊��?Fl��?�t?'��	����$�K�E�?J�j��O�3�%�b�:�#t	`�8P��u�����m�Sy7��Ց��f-z��`�"ٌ
}��x�>�a���`v�6�T����b���2������҆��޸�˂>Rf6#ǐw����/D�uIl� y�W�ǖg���S������#Yt18b��f�g �,��/�@���Vm<O{��2��[�"�c�k�%
�H�X���dL~���+��#d�.�Mf�����,/���u i�*����sE�WK;��!L�m��d�G*�~���M��@]���� �H_~Ģ@�;/�H�𐠇�U��I'v�L��oy�����h�bCcp�|�)c@b�Ɇ��׿����w��	79��{/��_�ߴ�t��$��ߝ9GH�� �W��H����|�zg�)���ԀIZ&ʪ-�*"�pl���k�ʅ�E.����**o<��0Ϟ�kp��B68��
�"qaZ���ֶW�W�,|��&[��M-<�c�A�\�`�U.��t���9ND�q���9I�m���q����Pv����]æM�n��
�'�FQ�k�!%e]q�͜ry�-��(m�	9�*��}&�V
�s���1�%Vrk;���j�]vO��Ӛ�����y��js�"7&�Ͱ�U�oc��s���D,�>��C��qt�9�CV�C� ��Ք�F�Ab�͆�ag��V@r1z���ȼ��W��VE�D��ͤ+x����>��qڦg��ݿS�;v�$+��4��؄���$���.�B�]9)#�)'��5QN�S�c��c$��j��IV���P��6������8[q6�S�w��)p�3!�
9��y0<���m�e��d1 ��� L̆96ſ1�n�"uX�Eۍ{�ܴ��N~�=e�+�@��1���w�߀�f*E�k�I%�[B%��((��o(=�X �V7�*�{�$��_�n9)�$8ժ)������i.�BuL��1>��]p2{>��3�y��^lM;8/�"�#�L&n�����͢k`�!����3v���觌��h:�z'�i�4ݝQ�����aбOW���D!f5�K49��^g�7��O��Y��Z��߆���Mb�g��i���\ќ�̓��[����?z��2�@���џ�<9�i��xe�T��Q.KFR������:�0�Z�ҽVN�L>�nl��"���z1�S�����?�X�������W��{��5f�ml��Α�*��A�<��l�P��e��Q4��x�3�����xzu�~���S@M*ro��Ϳ��56@�����p��\�k�z�x�� �^�O�{
2���������p�J>N�0��)ņT��qS�"�"�������\��-��́��Ѯ��<^ c��o��Ԇ
�}2X`Y�E�b��GF�������L]��ǥ��ӬG��?z�C�ђ�o�� �br�7�,�b��މ�Q�@J�6O6�����˄1b!G�7>��3��g
�ĵC~�v�1��m������aO�p�qd�ǩr�E/H�tfo!���1�їHp6T�_�v ��7���"�N�<(cE�6�L��~,I"�J"n��t��P��bY8�s{�M�=l0�/؍�_�ĹK�R@a�v�v`�h7z�I�co�=;�$~��(^� ��*+v}.d�5}�$ Eo���ǁ?���v�[[c���Yq�����P�)��R���\���d����V���|���`���k� ��h4�.6�`���'���$P Z���/�N	t�}�:?���P����΅J_���a�+z�K�w7YO0�`�_HyAy���8�	��;jH~:���\`�m\�_P1�Y�=�7~����O�j����:��ASc��	+�����q.F�0�w8,��tպ���������j��#*Եv�e`�����ce�P+ǡ��w��([���׎��=J��Tߚ����2{�WXv��nZ<��Z�O�;�~&�����r��������;��܉4�M�P�*K��4Μ�~B(��/�^�x z�H����:��>C��w�[�<>���5�79X'�H�`i}��%t�,�}�d�P�=�M��~��H�+����ǣp�t��ݚ�����:�j��z��2�9[���8l�>����Ԫ��-)G�z��L⪰�9�Nh�[�����gc��H�!�M*�@�d|��N.�R�<+l!�Q���T�ᔑ��?*��Vl���^���
O#�]���#��*�ȍuƣc|�Ǝ�9)�qJ����M����7���p�	��Qi�~N���VǇ��N��
6�衲5*�F�v4���l W�"�3������q���[� �Z�H>���U���A�x>�9[�d*����И�4���a&���'����%��8����dx�E*E�.^;�"�Ԑ���f��S��UC0� 莆��`4��@��)��p�礧^&\��(cf��o腟�?�]m�����>�X���`C:#U��,Ϡ��?�8놇��"�9_�u�;}��B;i\_R�m���ބ���V	��A���>N���m���?��l��$�u�Z���^�Dĺk�ɦ@k�������\򴆎w�)�%02g:ǂ=P���a=�L��T'n�(0�b� a���hTb�
ҔD{� ?w6H4��R��W[�gW@��T��߻��`k������~���b�CK&��Y� 3�pw��w�:�泃Z�V�Y�f�d��$�w�b�k�Ԋ���["W@����;�Aԙo&��iye�-$d,�|�ƍ��ՙ�C����MCwB��uB��'�Շ�|X�H���Q�!�IV"6"�&sS����w�^�n?j�?K��$�� ���brCk�%��_jA[�g�n���?���ԫ�1-,�E�Cs:���Ӭ:�a�'�4�S���
pMz�1۝C��a|��j�O�g���-N�a��¯��r���4���el�c۶�8�iD0GeC����M��������6SИ,�6Z���S�
ٛ+�	a�@�B�2�ҵw��"a�#�)�4����ފ5�V����1��{0���l�H�n� 2��S��-o�'���nR�y��Y��Q���רc�"��5��q-��ӆCQ�ˡ�4|%g�� ��d6� �߭:����*9O2�6��+ώ|?NUp�^|T��0����Vn����{r���ъ� hj���[�1@8����zU�S>;�s�l��
�M�U�$�nT�^�#SVm���N84���؇_$w)1 ,V���rU �^w��]�$��@ݷv�����`���<���O���0"/9���5n2�:Z�VMn��F�H�j�T����Mjt񱂋U� NЀT�4���r����E����g�ew��5�-X�
$+z���4�&�b�
�5)9�������+.L*j��P�Fm͆)�����2.!��� �$r%y]�2ϕ�D���B�yu�]�ac-��j���ž�>���>�Z7���3K��^fI��B9�\B��&�m�׋Mu���V�P�E]�X��4<˻���)Db�jӲ��1�o��|�8B�!c4��r\ѿ���QyEu���`�n������S�X�����r�[#p-$%��J���+��G�{l�vX����������r-��R������Ux16�(�[)�+�-��-%�ռ���VK9ƑLX&-`򟟒�p�cr)ࡖ�n�5l�>�t�6�׷L��|aS�Z�`�S����/��k��%�8�<��4xy'SO*�&�f��Ά�O���5�M޹d��o����Z�)C��>�d'5�A���p��az��t���'���a��1�4�Z�Ⱦ�-�b��k��t�oK�<���㽍�Q�4p��v���z�<BE3����2��BJf�l>�p{�C��K2���g�Y�o%��>D�}Uei�}�}�*�4�F��h�c��Z\���	0%�x�]��a*c4y�n����
s��Q��M�C5b?aԗ�k��x���yrG gEt�����r���@�\��������Z~�W(%Y�C�����j�·��%F4�$5���!gb�R� �z1��)����]���g>���^�ؾ0�f��+�T��ԑ������ƞ@>9�.�ȪZ��ڣT��ƥ�T�K�+��x��ڥ{~X���&�*�����B�^��u&�C	���r������e,��;�4����݋��"D!��Z��2G̑�#B0!�z�҇�88Y���}}Ę�(����l��׫E��Y�]3�Ǫb�{W���0E�kE���b̞�ej����	��#K�mY�Η�����o���+B����Y1�3����
��-`�#��3T��������m�����gD�6~��崻V=�k	R�� �R�]��p�+��Ta���U�|DE�ۡ�D���W3�_WѬ4��kϊ�ؾgJ�ɧl��4��1/��u�Ѐ�P�EG*�w��ۮ�u�'?��|��Ph��{�!>�ܮ�İ(��׉J���r/�R�8�,�����v� UCԽM���x�3����R���v��>�?��ٚ��y0]�����#/��/O�<p�5�0ȸ��J�]w�{�C?G�oO껻k��b��B�#o���/R���&S�&s���b�]��4��P�J�*�b��<0�;�U'���0�{b�Y���O��K��y�X�'`�JQ	�&6���K`��%N]��Tz.��Y�x)������ԺB�06�v+�2��7Sb�|�(�J���m�:{qn^*�k;�_5��O�xٿ��?�熭+�.�1��X��Qf����gٳdКf�(��'��]-�Ss��	�t�έw�?�c����7��"�Ў�dө��,��+�S�Μ$/i|Q�S�D�A���h���-)�������7-�$��ʢ��H.Q�('���b�>�׼H�@�!�]xeK�ɧ�ֆ���,�Z>�g�A�d�>���@�Iu�ʳ̕�_�k���Q��j��gY)lt
6����V���,Vxu\�޳�տ��/�y�fT�����`lJ����ɡ_5��F/!����.�V�,�[���՝ܡ�$o���D���@\��`�w����|x�H�`��q�]�D�h�$N(��Z	E'��Q�n�-*��;�G|��Du1qM��h�����m}�{�e�F�B��ޅ.?�zȦ�P!Z hВJ�R�&�
-8.H�kh-�XOp��G��`c�I{u�=F!���fS~��C����h�}�)�P�{"U�x�,lD�ړS`�/�[��~���?��q?������bp��yz]ś��-�?��f�E�3���VxU���-ӈ'�w$��(u�5GH������ߵh�ɐ0�7��iC|�T�Vhm��A���R�J)�-���wS����������L�m�ͽ�?<�u�]���81�!�+�$�����=m[��h(���v���Q��4VPbN)�i11q×�a٪�'ru�oh�ݞ�"=Ѷ�"�����T)b(�����}@�Z��qwӿ�X��V���=�.��Sܽ�=�߼�UXq�W��?�M� Y�qӔ]�6��&�s:�[�b�i�5�	[ݧ���(��Ap'E����ql��̉��O0fb*��t�Fŀ�$�A�}ߏ+�8���M��Ҫ�����HO}�fc3�*u�ܓhࣿB��]����]��o��W2�ܖ�S%`8Y=�S�%�&	�[��Km�;GM�"��zj�$���NA{'��~.�o�A��M9'��&Do���Je�Xv)/6����sY�W� �G]hWU��%��P�kF��6f�0O��4e��B����%3I���4�yf���}�
g����Z��ٓƹHvuYᑪ6u�Q�`7=Z���ÉWj��^����s���7�+�{]G u	)� ��|�-�|��%d����x�;�0�Eջ��YT�1W򻞊�%�N馗#|�LLq�1�B��?�+}��$R�1R,�ypA#:Ɉ�2h��\�ś�Z��x�ЀJ|珂n� X����[ �õ��6�#�{%�����:*\�F��)��J\�z��%�M��K]�H�
�Ol'���*�)����E2��8��!Sp�щ�|5���D���&��>q���@�T Y��v�V�#�al�E��ԍH�R8�D�wI�S�4Z�D�6՞�#z��a	@[���U���=&hNO+@��o�Dނ �mbݜ�'ڱ
py�R�A��P�4k/)���-��F��#�@�!�d�#�6Zp#�-}9� t��C%��j��1�v�j�2�Wq�I2�1�8����q>)8�q���u�`�+I@�7��S�&�2�l	�)�L�^e�ѹs��#��&QV�����&5]�Gi�-n�`�%�͛\/��x��Asv�*Nh�Цс
�;���*@�M�$��80zNJݛi��l[�@�'\�6�AB{��z82YO
�ap��
vr���ZA �����V�b��J1A�H����נʗF`Z�f��V�ɑ��/ nog�"7��cH)�e���FU�����&۔��Q�߼�[�)�����B�'�@V�ѝ�G�^�!dd���X"%+� �j`�3�#7e��(P�#�m��N�
{$��ą�s�;�[�֊��
��$Յ�R�q�0�ڨvD���� �غJ�1Ռ�X�8�&1��G}v١�4v(��]o<��!+Mg��ɗXu{�L4�
�F��I�A�>���P2㸁"��2D$���v�*�h'�E��Âs\K�3��e���Dzg�o�֞i8xy��t���L��
�l��!vB*�E�q��0����nw�! ,4��s���l�C����ۮ�Vol_s����z��.,�C����p�t��=��Y6��
�ؾ��8)v:�J}-ȳto�bsӉ=������ƾ�tY�>�=���3l��~�xp�aƂ�� �)���ڈ瑠8����*�'����)�q� AX�˂���CΈ�qm�u�W~��Z�AM��f�hFOm������o�P>㋣�i��ze�^*�H�2����f~W�.��=r٭��Q�7���Z�Fx�.���gUĶ`��v&�?��Q��RCvζF/fд``�v�؍%�I���`�n���	1X܌�X,?��D������p���*��%4�8Ż�=���GZ�4LwԾ`SA�	�)�`K�*���;v�K����@ ��6a�@m+a%�2���4q��ԝN� =S5�VM������fm�v�9���/
V�Y��"Bn�E��ch�<� ��YA�;���%�!�f���'�L�x*�
4s~�4���>iW�
���6MC�+�'Z�w��\ҥ������0���A�RI(���Q"Yr����������hHr�5�e;��0�&��q%�� �S֪��P;U��"~z�R�~9��'Rj��jg`��JM��!joմ#U8�������u@2��Y_\�[���)�慫ϴTt0�-��D�-SP�}3���c47�X?�滌Ŝ�ׯ1� %Q�"�H�)���};�"�M��LK������k������
I��f�q\]��^X'�C��:�q�$��m��d�)�g`�Bʒ�I������U�����Bۍ�Ô��-�L���c�sߡ3Z���s㤞b�@��G�b��տ��e��33yn��ճ������+U��p���~�8�Ca����BGjby��� :��j}0�Ge?�9��r>����?I�C��٘�}A��ī��E�T��h�Ir��6���:�Ӳ�����?T�]�oY��v3'�g�DXF��+w���������vJ7fOZ�P7R�����oM�τj�N�h�s���р����xJ�d(R�O9o�g��_���=������O�9k��w9h�! ⊕A�w�1��y
Ti�9�I�ebĕ�a"_}z�m�Ի��r��@�i�~�.^{�Rx���^s�vi3,j \�t����y��M4��ׄ����`�fp0J`R����혬1L`�|�āE�	:h|�6��z�7�;q���P!y�B��Zdu@ࣿ����!f�l};/�@tJ��<;�D��^��-��s����VQp$Þ��[*���G6�|��
�^/�B� ���;T�و���4��ٝ�X,�LʜS-�|+��7d��6���g�c�Rm������ �k,l<�_M Yé��N�OC�} �"��'l'�CWKb�<�)�L�h��j�wGM�&e� ���V^eQ#ri����Č�݀.�� qޕ@�jK|q�X0	6��ƨ�&�JG�	(�� ���kS�)D�_t�_M�7>��yrc��V���u�Io��	Y���~3�t���46�����fn��r�E[��	{gk2m�R�;j<�ͱ\��О.\�:Ҁ"j3�g+��x���3��$R;��;:�;��y����N��#��<��_�5�ָ���ې-���Z��ж����do�K��+9���`/\����y�GA*m�Q��Fۭ���#���V�I������g�
��[kV�'<�W��b�aq�.�}R���ߦ� �He�ˎ|���^6+�s�4^�#�=o������{�Wl���,��I�'pu�A��s��˃�U瞾���A�����EF��x���v��7�K�e0��&Y�]��O�*a叆cب��є
�'d�92���_��O�����xǋ)�?<�s��I�E~˦2��T�K����2���	�L@o��?=_�Ư*<�V��k����OJ�	��_M���j��fő&�W
�D��K2q�_2N!O�BÊ�,�		s�(1�D��8�7��gn���8~�V���J�rbn����U�Lܢ��KY���r/qD֖�T���~L�@Ͷ��A�$�C���;|�����9y�s$1���]~��^ˢ3�QD���м��V�NϯE����uU��?ڱ�A=�^O���C=���h�@�9��+�UX+�V��o�eG��4I�����@~�� e]j���/(z;���O\UF������?"t�����\��(�ѣ��k�i=p���'���᰻�k[�3E=o��Y}m�Z{�t���:d��C���Tfe�a�;-�P�ٗ�J4�]�$�E|m�ͽ�#��aHϠ�h�ѵ�-��=�5)KV�x��g��0���@�.7򓞮�ی-b]�-rv1?PE=����I ��c�Bc_InDեC�=�)I`��X&/���ay�l���`5�7q6m�'5�;DњŁ�#̒
����*s�ؗ��L���.�#���ǣ����9��o$�%*�.�
I����ّH��J�A���2���y(�2��=�{�z^����Ss���l��&�|:Q�cx�3�;2w��Օ3�|���3��Aa��ݛ���腎������`C���� y�T�F�n�t=ւ+	ЏBF���	���6Fi5�^Ĳ&�~�jS��a,��^����p��N�0�`yx��]>��o�)�^�a���@�����t��Q&������׾����+�;�B���OG����]5c.��zyAx��P�l�Oߗ� {��L��q9Q~���Һ4IXlkbΩ���N�mݺa^�|t��tE4��.w]��0�Y�$%0]{Yl�=�5�R"YZ�l��,��(�[t���]��p�?Z���̺A��{�	W(����p�y��<� �x��g`A�p�v<�]%�MɵA�ix1Y�h�
SXR���Q�P����#� �Чj�K��ΆRN^-�_Wp*�L�6wi�	~yz��do����?C�X�r�X`�)�9�"࢏�����fPYٯn�X�� �'ÿ�[�X�F!����cQ<��N��~�~�@gN ��-��A�үj���d�^���(^%q,�Ґ�ī}
\X&�g��RO�g���@������	Y� QӃ?�_��l�~ً�.��)�	��}�h�I

+p�%�RE�b^�w��3+Ο�r�7�v
v���̓��f�űE��9�>A��=���/U��CJ��}���/��8U?g~����Ҕ�m�n����: 3��V����������R� Y�߽��/�D"�'7]��2м5�1�|��|���_��i��f(U���M`�["��/��73�m������&�Z6��ѩ��*GZ/�y,����/ϴK�n�����
����%߈��������]�B_��ѼU~9́>�����!��\������#��(i�,N����o]\���|�4��Qɢ����m�Zt-�dSKIo�-V�[C�si�r�@�D��!���ɹ��Nڼ�@6�ȱ���S§�q,AV-�n/�@�/��}�^����^ j��S����?6���1I�#e��*, ,�J3�諎q���Ř-쇤����?�vo�|f�'z� .���V\����X�T��x��s�?�'�+0��hJ�I�uq�d
�@�A��1I*�I/ RW2��';.V�w����w�hG�S�N�d]��x �a�S��yH��|�0��(�cN����Gs��/��׊���g��J��MI���۱��������7�ŝ�:�/ '��_��J�x��=�t��U�[cP�b+ݪn@p-%0��y�Z�&(ꀒ;�6��o����^`��s�K��{��fS]�gB���Y�խ�g�_:8TH5��Ƶ1*z����x�'p�~�,�=�v���e+u���=޸m����N��1�W2'n'�S�xF G�h�H7�j�"��2��`P5�7k[�gP���_����G�������$3�̼�c+��)�Og����wgLڊ���{&Ʒ�֫<z��)���A������R�v�Iޛ��7"+	ہ���ß��j%�I+I�d����Kv�_߈�J���#Jz~!?��xY��S�dȘ�3��r�6]���m�wQ|e1̸)T4iɄ�S��\�N 66-	Y��}�I��Ї�)�|�1�&����܂-G���s��-����/�L�T�p�L�G`	�(g6���f�������*
W���6A����������K�U�����ʨI�au�C�͞��~�c����t��a��C#�t������%���$"�d@�¶�v�i���=�cD<*~���j���@d5s�O�M�p�C�B(��c<SNd�09f�R�b؍�N�	ƕb�r�3��o���@�'�f���s����2*;C�o�U��Y��������V2Lrtwo�9��d����"�#���ǎ��h\�Aݮ�{#�-q��������Cm,-��;���b��>ꌂ�P�����*�D4�
�2y����P�9`1U�'��<��Z�:;��DDO`Gv��$��",�V�t�)�[]^�b%{��ŕ�?ݯ��H$�>=a�+f���)Gs��H�������;��"�%��  � E��5�pJ��r��rh�9��F+/J�j�7���j{3���>�� �H;C_���e ���
�Ek5��Sĥ��U:�R��jwټ'������	�����5~
��ik|��)?,.�R��}��-I[�B���H�tR`iKdp�ޝ�k�\ �P�a	��4����|�#�%q%���u�A�
��@Ki'߅��o�e��2Q�K�[ܤn$|������m���X=�@f�؎{ς (3QӼ �����o�z�I�����q=���P3��4�G�x�-q�@�'�J��n�B=��n����m��j��S��JA����BO�E0s�3���9�h��PM���>��,���WU�#�	�\#��)i�E+���������t֚&����kg�1�����L�<�3%o:[���!��;� ���+v]�h��m�37=JNF��-:!����Z-�֯yȻ�h_�QMKz���Ot�'H $����9$��CO���=���w4m��?A���q�t$�@���Ev=����N!K[�L��)�@!m
V6l���2{d��`^�r����/7ipJ����̇���R�4��ߢjX̋eᖋ�-��z��3E�/��h-3��#Ov��a��W�O��s.la����
��r19I���ⲏG�/�
Y*��X-m �O ���'.O.8��z��m.q�m��,Zb�+�y�۬e�w�g��N�e�F�}�W:M�Ix����=��OE�D�)�kgf��D������璘�G`2�M0_D��$�c���1�&��Aܬ�(���~n⢣�	Oˢ����=o�G�W5�K�*���ϼ�L{�5�

��`Ϊ_F|�Fw~(�zqc���_y@x�����/ ^��i�ɞӬyt�,e��⛳��(?��i�����\�j��h�y2<�>��6"�i��<'k蝹���`����f~�'��v�ܐ
ݻ*�yF�p�j� �zϞ0�uݞ��7or}Z�c$���x;�<솑>1ј �XD��ϩj�M��^�RK���8��G�DR\�4}N���g������}���KO�y�Oi��T{�L3c!�`��È�Q����{�
�ޤp��@���15�9�/k�UFn�;���H%�o|4���I%�+$���Y�~��b�eG	 \}�����<1j"�Y����������H��J�k�>�=�QӤχ�[rϔp���ӯw��o1Y�!��������&�w��.�,6f�=�C���f~�Q�X��>�d�ow���	�L�T[uzs��ꖉ�lOz��K�3d 9�xGX^줷��/(TZ�/CF��Yoa<t���#�b��%3NR �)�
L�Ǖ-����\�Q��@��{;�=���>E�1�g�}n��}0ĸ�b�PS�(� Gݲ��j)�V���q��"&k������e�
�}VE�tѶz��R�`F�p��Y�}�RU�P���ۯ��.Ob;`��g]k7$�9��j��/�e�<�i�� mUi�dۃ>z��$zT5��OM���i�7�\�����K[�y��SK��qҺaEXů��r�"�B���̤g����{��n�bˊJ�$�
��x/;j�h�Cl�FM������������g��Q$�h��02���D`���0��@���B����������-p����<� �b4<�K�Cd.�.�)��!����r�;���F��Dui���â4�x-"S\��(C�)RCQ�c�-��;݋g�}#V#�!R��6�Йvp*ߖ߆�_b����X&�Ƨ[r �aW��j��N���¹<֣~�5���oß����UAMqG�S�w��f�37��R�ˬ\S,_w�V��ḕ��YCNw�x��KG�v�z}�H�����X�9���������JR�#W*J����;)0��v�DbᩂbLꭡr�C�7�.-"�E�7�ڻ'����1$�~}$t~�;v�_�+���/�*�b�u�o-�#"zBȅ)�mk�5/0�R�2����\��6��=�)Ѯ��c���jK�"�(�mũ�>[9�����n,4�F08����,~�� �&=<�j񺇳�e>̠;L�j5ao����?{&e�z�(�Ɋ��n�7�]2��UP��n,ַ �[����/a� j(�秅��1�f��G����rjd��j��)��R>�4�P��#��<D
 �C{`��	V\Չ��ϟ��rjF�f�����9�S�2��!�K-��DXjGx\�2n���f��)�(S��upo���*��2-�5oZ�n~�D��}$�q�N�7Lˊ8K��'$H���Gaԓv��(�X��yI���e~��afnj�|ѿ
�W�ʧh2����,Ӿʋl�K�iS��y���,q�},pj��dc+`qQ�|�D��8a�u߱a�7!�=�҉|]�<3^�4� .R�mb��Gj��"�̐�3��5��������P�N����P�ݑ������'��	!{A��s�����:4̮�w�-�R(O��0|�� ��..>�h�	:����a���Z �Kx���7���T����N<��_6ȝ0[�,��{�p���2o�����!}[��;`DQ)Z@�Ցtے������^GֺXB8I��M��w�G8�<�x ��f�ԝ{�
�%�4�mQ��4��6�5��ӽ�k�R�C��S�,��s��e���!(��z[%��fv��"���֐�cU�����*��җ�=B�{���K��Y#p��,7�;��y9m��^q��K�Ɏ���\�-F.���2�D��7��ܰt�9'�O�E��=*��V8	.�?��3��n3����d���2b������P����h���	�rG���A�q��;����j�P�G��	#�S˙�HIor��!�6�qU��_�N�����	�����[�<ȅz�.�^���"�K��l��1�#�Y:���j��mA1E���	�.N-�%yE��D���j�[A�;���YJX�l�m��2'�x��-�z�����|֠�il��ѵI��y8b&�/�a[�`����2��>�$$͵������I���at��D�ي�P���̷9�mj��^,�=�78'��?��=�BO#ٟ�N����,U��,�d�W8�n
;��R�֟@X�	Z��ұ���5z�ˏB�����i���`&c֊~���-�F��W�U��z˖J��B?4W~�(M:=Z�o�p_��J������u��$r��Q����<�D��R�j��aţ��ޟSf�T�nȶ�-�q���!���M����pq֒ү�Ӛ�tvHp-�t�	z�8�BN#�rW�7���񻭿��ȭS���
t�=5��x]F±��fN��P'�[��i�=�������cM�K%�&��7mc'��]<=[MID��2��{�3���~�E�`8���1cj����I����/�Q��J+�i��:����0�͏�
Y��~��P)�Z6.��m�Da#�|s�6��^$���GaɊ�92;9�<xQ���wT-�evN�_{C��#|�X��tFNE��\�n��{��g]}��/j踝��M1d}4<'Y8�<cZ�r8E��)��]z6b��Yf�S2�o����\AM�|�Cb��j �iʜ-� ��,��6D\�6:nܟ-���ҩ�@���C��6W����[a�w�����e�(\���M���������$Zw���Q6���2���خ�5g��o\������%Hy�}l���G<�be@��	d��k"}����{�>�{���'�1��d)A��+�����3 �N�ݭW�*x胗�ܬ��	g||����iE�����48Bb���
���L� N��+��>ouVr!�zS
i��@ Ɉ-�H�j\� (5�]���P�����$�4V�������������{[4��$j"�0�����9�G�j3��I�)m�c�Yd0��m�/�d#%��|�8iJ/����$���@��;��#��{�R�m\
Yl-Ah#h�f����k3#�7$��%>udlԃ�E6�8�U\���_���BX�މ�E)�T�|�Q�kFl�+�4�Nu�^4�Ӗ���|H����_�K�gUL ;���x���4nq)I'Z�N��H���c%�0�-���;�I $S*P�� �)�t'��A4k��4;e���(ؐ�D*B-d�D�
��ġ�*���ְ�L�
�T�J�O~�,�d{�mX.QB>>�cC
�˫CW%J����a�6��!�=J�����H�n��ߜ+;��4�"+��'��83�|$a�l��`�^����[2%x�ͧ��]��0wm��X�-.r���	%y��S�Y�����q�"������,@n ��ck���J�����Q`�aQ6�۶ �I�h{d�����Q/�����䣛q[}��⏊5��Sv�a��ea�%��^.X�+bE�e�[�B�$���G��g��5ۮR r����ȳ_�w��7���
<����|_�B+ߵ�;*H����W�}YM����j������;r�C]�D̎G�Sf�RG��������P�Y_N�s��o�M4���L��Q嘌e ��b4���Y�S8R"�&�T���s9h�Q1�brr�sUaL�0�6��Zg�x5-�O\��I�3�X�Z+��J^1i1f�}6y�I�oyrh ��z~%Z��Ep9Vb�r�8Q?#���"���3(UH��bW�F|�k��qc�_�b�ےx�c@�q9�Zz�y?��	�5�I$qq�J	fŐj�N��ƥ��tO=����'��TMBW,��oZ��6G�_�7�Q�a�����0q��M�vC�����?�;�D�\�v�pۿ+��l�� *��
�T���ؼt7��(bD�^������D�4�����ǳ��4b4������E��������s�J�VF�?V�m��I�.!����-	Wo�ު���$��?�|y%�kz1r������z��3<�)�<'˄�l�#p�zv�Vтp;�k43�wφ��4rb^E9�`���>�Ί����d����{�j/�7�nw�K��5HQ��{�!^k
���R��@�1�>�!��3n&�Jn�l��I[�o\�l���c9�qkcε�]f�\�Gq=U~e��$n�t��}�yY��<�b+��x��M�P�Mܹz��L��͡K#;�eisfC���֖͆X���ڟ�^�_cb���=f��Y��� Kp�Af��t��W�h�܇D2s/0�,�cw��,FM��Ԯb].�yh��~��V�>��+��B��tb�����o�8v�>�${�����鷇/v���ud����'�n� e���钒����PEvdb ����7F�F���b���K#����*N$��G�c�������<;:�p��U2C[LBF�x�"0eݗ�#���jX:WX�����VQT0��ev�ۿɨr���M6����.�g�d�~��{�,T���t�\�x����P"�A�:��h�?̖��ļ�}��W��B����º9-�Ó�������S	���0�K��Z��F68Q����	�����x��ȁp�p�uΝ�M��d�zZ�K	@�5����������ci�9�`�;h��q�4�w�F��#�DM���x��q=�� �Ӕ��6Q�h����4��d�0 ���v_�����Wӳon�j����i�6����í=�,O����70-��܏f�ߢ�V��[�	`��K�d,�w��ʃ&���OT=��[�a#�ߗi��~}1m��ߙ��Z�h�%�-VH�Yy�>���+�wkSaa�����l[�����G����`���;y���{H,�Tv�����T����G�y�>��i���-��&� {�>�l�n��;������Y@�A�OÄH�OB�(!G|��J���f�np�f��>ֳ�_>-���:�k�7l��:�)~&�����aR�7v�=�AW�q�|;nY��=�4�/��P[]��}�4'�N�[Q��?�>�)��R駐��'gP�KPHK"ew:�w8�A�/Đx�^���x�)QԴ�	�H�(F���]��J��שH�X �E��_�/�є%�O�:�������I(��%8�@ݫ!�9;�"'���,��w|����ٽ���;���0f��<.W�Ҧ����W��}�����43Gi�W�*T��|��F��l��$��x�����r(�GuvNtSwv��Rk�[��X���*���8^�d�9C�9�5�p��N����ٶ�)��6��W�N&�'��nD� E�;k}�%Sٟ����J�C?{��p�aIi���Ѐ��[ ��5Ŕp}�ZE�|ŵ�0��lR,�:�qO�����ʊ��0�7	t�:�C�H^��A*y>�����S*�ӯ���<����x�r��jf��w��*@b�鴼rNyV��n�8@��2���� �^�����m�%�s~���G ���8�lIc=:^!]2[��t�GrF��wa�df]}���q4Y��� �?�Ȧ����x@�\p]mh�\}\F�&��߳K�a9�pډ���6�6>����J@G�#``e�_v�801�tO=���ȓ���뾔sS<?E&/���C��XϽ�W�+�V��{\`v;�� �I���-{���ޝ=��/zs��)��>�~� &x����2W�N�~=���7�s`�z�g���*�`"��ya���\�a��\�C~�L�kK��G+�X�#Hj.�����k��X���U�gIC�P��+���P�ۊvT���A94�Q�0�;.�w��i��"	f!�TG%4��@f���_�ط@�}y���!0!`X�0�J�2�a�9�n�7@A�B`AD��V��*-�@4�x�̪�8�7�P�mŠ�;�f����s ���a��H8w:��`ϓ1��d����B�Ƨk���� �2��4E�p%�\�<�钇�H���ὢGh��-y\��N��ۨ�q�C���]CX"豂�.��;�}~o��Z@8�p��*��N��f/M��M0���������|�Mu&�\aU��#��d�jM{}�ք�j+ʝ�!l���@�i�_K���& �U��U�wp��Z��0W����R�ui��T@URcg���E:�
܇"��vJ�E�xa���Ҟ�g��Vܻ�N�wV{��)�q5&�,)HV�{�z��ʒ /-!}g"g�ML�6��
��H���fk;���s�� :Kj./DַEk� �/��R$���f�`l��k��UBs���[�H��~�ЊUc���������y�/�>��'d�)�/b������~�?N� ����6�!\�Q_�co�CB0��}ی�c�(�(c�Z����0;eĞz���셑z�T�I�Zh�����΍N	������(�ȗEy�kP!��k�͂�ݴ�6�v3��Q��g(�>��ѫ�C��j��J����V���/A^�MV~��0��'S����e�}�C���]uJ��M��hk42[�W2�ھ����΃�$"�(+����VL8�Δ^�~�ˠ�������ۓ����A����m*��$���	��x:d��; m�GP�p�G3��;gh��A�B i�?:u:��C����p0�#�.H��|�c��^f>�}�N��Сp�i���I��h�9�!�u)hx�R��B_`$��4^�����"P�]���?N��a���7!T�+̞l��B�"��X]*�X�q�uq����5 ^�g�Em|�xW�5$�r�DSB#qهC��t��KC����=j��N��!�&�p�i0��a�]��[qoF���K�)�u���܍�u���o̒?c$L?�u���������X�V�����T�;��\tvǣ� �#�8�t�=
*���_w���:C��-~��yo@ɳ6�'���Ŕ�q�ᄉ����j�	�TNC�^6|�o[?#�-��kNpm�1�'���R4AZ��ng�I+����"�H'8�ʅ�����uM��b��KŞ��gl��и��q�k>^�CME���Spc�R�B)e�"��Ck������+Va�{<���U��9l9ďh����XB�V���Ŝп��P�z��� Kv����B����[*|՜U,�Q@2��(���2k�ݼ�����0�O��g�6ni��	�Z�D�jyJ���������~�*D{�ŝ!n�6�J�Q����a��xD�~<�����c��kzUw��_@W���{J��v�	��K�F�1�&���@����b%�?�mēj�Ca�B�v�N�u�!�#��}���{el��6������)�!�9t������e>�T����1���W��D���V�z5��)  �> ��-��ca�?��^^�!�G�\d�B)���2��YR*����
%��Pa���@R����V�`�U��h��Q���	6/!σ3�m�ſ��Vn���9�c�d�Te����:��ϒ��A0�����F�]��Pg�|����T����禎��~TK��6J���T�_ �x;��xt��O�.�tɡ>�m9�Xe�������&7��ž˽��^D���=�?RY���4g���\C����ɽ�s����l�s�f�).�ak�kЎ�'v���� U�)7�A�;��GY2�<5g� ��L��L����}Lv�\J+�x�ߙf��*�1N2��j�a� �4��Q�@��}�X �r
ch�����vO���2��b���x͆#�c�z�ޕ߃6F�}/�?O[$z���k�H��~��	2�OԾw�,�E�� ��Y�Aa�3��
��"�:^{��(tK��b��g��1)������u��*C�gte]+S=J~N<���fʕD����R�åT��i��A�j<]��ݑ!4X9s�s^�*�5�O�c�vj��6_��A���86-�RQ�V-A��.�#�J��D�*K��'/��<�2��Ā� m���^�[Ȏ�!�=Z���rxe7u��ʾD05#��h�!�H�7'��fP��k�w{�#Ƚ�N"�����R�a�~$�F�C#��h�M��	3E��P㡝t1��8�z��ի�SL�L|���<��[�<��|��Ε�iQ�����-�����~�Oq�c?�;q2���Vr4�>����mTV+Lrt;}� A��"֨9�~�k:�u��+����Z��ƧФI���KS�RVĹb�J�@�U��Ǹ4��.��--���u�3|}WH�"&JWwy�z~����U�r ���\���i�;ճ:3� QdPh}�L#"0��:��Ѭ�s�]0�G��Bڞ��C&�v=����"�Vg���Ш�ݰ��`����
�k��h�5�"�Q��y�,��Q|ӫ�?~|:�B�g1<�}��?���$~ۿ�R��U6�_̤��D$X��ތ�q��2v9�h�p���T��6*-�D'��nи�[���8,lק�'������9����}�K<3�}.�t "�G�Q 瑿�������Erc�z������|hn8OD�"V'A��7՞��z�� 4LOp�}m�t�8%+�Q�h���&"�+T�: e��H�%���32���P��H�XBͩ�����\�j�-{����s�.���Jdi�oB�ĉ,D�Rhr�{u��ʵ�Βs��o&�� �ڇ~�	Sx�:�MzQq3&q���%|�-�Ĭ"��j�4cG�#s92��:[��o��sb�7��9h�����)_��K���9�ː��]�k<+���98-Q�5EX��8i����n����TM�Aέ]��؛e��`M}<N���A�p�Pw�~Ơ��Ah4@3φݖ9<�_f1�XktK�Єq�:�U�@���l�@�����5&��ه��Ux�芛S-5�+y�k���o���ywW��۝��@TW�Z.��E��Xv��x�@=�:��QSR�=Q�����˗FMS�&�R/��,V������
�ӂ�����'���8x:�B�nr���}`r=� �Ǣ��K�Iׇ�4|��ǹE�r��@�*���;[R4MB��s�Y`�w\Cpl7����ۚ�NP�pҎ��"?.�	���2��,H�[k"��V����@`���*@[��"2�Ev	r��JW)��YRG���D,I터=�_#�9��ƘGJ��?�%�m8��ܰ���w��I���_�\fk�U��}�.�HV��cqZP��t�7g.�Mf	�H������� ����d��e��شx$P����67���(�J!B,+y�SN�a�5@�|�iQ_FȌ[0�-�1]Z}���Ja�~u��-N���_�BT>�2�4�H߆l���k�!Gٝ���h���e�\��Ɵ��J����g0��ܘ�vR��d(Y�YLkC��b?hżX;�	�E��ёL$�Dp�?r�8.
V���8�4�d��,�*c2�����Ob9�ރ�#�}�$R�/��D�]�S����'��V�~~� I?Xi+�b������A�r��Y#�J����6qd`�:�V��L�b2�.�YQ�6�e�<��s1h�]�g��wF����h�[�y�蹚��TCų�9�*/�?Li�S�u{y�6�զ]���z���{�X}�
JJ� U���[ԕi���u���.�<�����>�>IP�|�ι�(���l;�%Q`��4���x��v'l����5T��M�43qu*Dk�wX:k{Ye�WG�{*��|�:�5��C�0���mX�)����G�\T�˫��z�{�@��ö�4��;�/쥵�Q�Y�,6P�,�A��F0�W�-f�����n���1����Py"�;1�l��ݵ'q��<��a���̹�gs�����l���x�Ԍ�O(�/35����N&;�_�惍�2@���y	�]�o��&�BQc�x<y [��\ޚ�<-������&��:��~�U���uJ�X���I���:����p��"~{��I��u��!�+�D�����Z��Hx;����Z}����J>m�\�B��k�2�*(NE�<�ocw���i�n�~�a�bB�7m��  ��-��W@��?�1W�혗����G�a^kzgCZe
�;#�d
GM�f�7I����.)X���y�$�Y��wQN���7��)�^��چ��ni��	��g��Zm<����Y��s��{�/2m����-��Ch|�=I��ɸ���;1\`��%ϒ	�9 ����w�����P�7,@����u$��Xɕ�F	��3�ż�i�3r3��Îys�q�+a�l�4����,M}���-����Ƙ6(W����䴓��^�*�#���HV3ք ų�z��uiګ� >��#lY�nFt��Z����L��80+�������|θ��RmS?�W&��/��3M�l}�S���.�1�dB=�+
��]j��A/�ژv1 �� ����N� LO3�~a4��-��'���&t^�GE�48��麦k]ͪӤ�rK0a�߈�<c��$����h͊G�-��6��jK��6{���0W��|YK����N�t�3CK0.W� �-aRǩ��=�c���UN�^��d@���&e"�����e ��,)�Ɓ$c7\���@.']v �,T�m2#�J��5��G�q,��/
�ꍉ���z�`�Q��5$pת�c(�H;��"QA6$Q6L�d��o͎��nF����<Ճ=}hg�{� Y�n��@ʰ�����)��g�d!a�vNG�W7|?�	v?���_�[���M��f��Ki~&:��k��oI��T�Y_�d�����I��[u@��|w&�2�ui�5�l��K�`���!���*e����)Yvo���08u�o�����Y�1f�X���T)�T��c�۽��##鶧̎C�,�L4��V�@�������^���ml<�\�y����Z�#|��fa[�:_�0�_	H����߿'@J��l��owIaH�@�!�bQ�p����4Y�-�p6�Դ���76����uM�6����e��J]N��L1~z ��+ )^�z�k������ly��{p�
�(�j��nk��`�Yȟ������m�U�m����䶨װBZ��.��B��h��X�`�R�pU�u�רK���MN�(�� Y�8�c�Kj�� ���F6��T`"�����QdS�5E�w|/s%&��l&;�;���ګL�����J�^�f@��h�x=$?�'x�[�"����e@œz�vY�@	�#�Y`5���I��p2wҁ-�B�����C�I�Ƞ�����'G�k�Ǜp�`.�Cw�o,���p����M����!�*��F��`T�XDP��y���wrL�L:�y����~�P��R$e?�[�$�6���j��R�%�R/k/n�jw�,W�J�C�ܠ��Q��Fظ��qm�+ I�q���LuXbx �(ɿ�2��K��� E�CL�� ��F�����L jsc��)+;��'=�/*ef{{.4�D6�	������+�<x�>6���
ȫ����_�GS%�B��Hִ�-��`��u�����ТBU;��ը\��`�̞�{ܵ0Fes�X�]5����ϋ�L�QZ���dK���t����_��Y�IRK�44�$��&!@�e�9H1jU��SC
,�����B@\�@T�=؉�?��Tc��_g�M&Ͽ�K' �_�X��|Z���\��%��9���zga�Ta�?P�о��=�13��ߚĦ��C����FN�s+�X���P�J'+����AI~�SZ�N���i>����S $�D��O!Gxlz��D&JL٠���;��X'��,�9��2��Xi�c��w&4�[v�B�-<�6�z��D�.�:8^{q��ڛ��Nkq�sBЖ0�����z��r�
�(��Et'��C>(>���l技�3�ik�9���HWD�r�>�o�ÜV�k������(�eQ~H�W�N�r�B@w�m�^���G^wޯ@�h�ؿ�U�(�.�蹰ɲ�Y'�å�3M�~]�����
==��<-��E��;Q����>��=0�ҹ;�d�B�`kR5:yOi�Ql�i�	-���zik�ek<d}�02%U*�N�~j}}�k昔p�V�Û�v[��6X�U�)4�	9�P��a�VORy�X6�)K�n{�.$�:�'�;ٜ,�R��������	��5!z&���>2'�Ta��EHe�>V�3u��ʎ*`����<�ͨ�����^�ӰF$�]�$�EǱe-U�z}�,��iW+D�b�g��1�g��WRe�K���2�D� .��0Dѹ&�c��b�4]X�dd���;RQ�z/���w�*�z��:�2\�i��/Q�+.�*��Y}1���k	�|EG_���V�=V����29�o:����*�m��
f��Oo�#�'��N2��7��~�;{�£n�P�(Z*�L�I�\���Gs�:���
������j�vܖSȆ�G�g�sлX�3���	g�j���0�Xؕ��1,��&x w��\���k���Ƚ!��j����*�t=>4}�OV����X  ^{�ׯ�F���#|Y��"��y+}��
�g�ٛA�9�\�#�9�xkI[Z�!H>Q6);�?��(����:�Y&�[c��$G
yn�K��뀺�<�ş��u�vo���)k㈆����̊��mn���J��G�%*S$��U�����҃�|�+7҆��4�2�ġ� �F���?�w�ODrs�3#d&7(]�0�(|��D�k{[,��[u-}1���\Zؔ�k.pZ�}�y��{(��~����C^�@w�L�)�8;�>�, �m�.�3�^�ZH��(��Ò�HO�:�Ti'Дi��Æ� ����Ƞ���[W�ij�F�d��ZD�Y��K"s���5z[�s"q
�yK,��E�������*r�;['�5Ʈ�й��s���2x#܆q_F���!H�)N&����JB�����m�؋م��i��:iھ��DZĞ��㨟��Cl���B��~9,��pM���J5�b�87E!�{D�s��iɶ�~����^��Z+�O��4"��WL{)	9�-����K_�9���̌�dq�a^ �\=�ƾ��kk�B�k��Ye7b�^��`�-9�S�98���QnF��^�[�XWIC:D�	�w���pR��x�\'%�Q��d�112��l�F鉭-T-vGg;@���3N��k�\�	Eh��V����ENs��h��4h�r�	����ʯۛ��)!��5��$Y���d��焠���\�mgf.waʀ�5��ݼ�"LE*�q�~7��E=o0�{
!���ѥ���(�r,��X T�ֿ� �߀+��>_����sP0�2�c׮�ک�T�B��N��?��ب�ns�qOW����%�МѮh�[U�����I&�!=�.6�cG������<���
^��DF��Rt�̒��@D͒���m]Pڧ�r���+�z�"O*#y�|���LV)Ԍ�Z�
!/E��֮�~��
2��'M4W"$��	���2�w�ڏ��";���_�$;��iQ�/,u�6^Aj�ARP>�5y�EW��ؿۚ���X�On�W����)��u�������@��\y����
�Eᝨ$��o*jP=��.��8���0��QY�Q�@��|k��5YP�F��O��!��ÒUN�]�c�O�w�p�CJ�T��;[��zj/����4�e'$ʾe�:��4U��c�lyP�z��d�Ǩ��U��b�-�x�Sʢ�U@�(����u������PG�h���1��ߕ�N[������qFi!� {ȿF
�kI�$�a4DN#��]|`Wu�"��:����
J��s�|&��kм�o�X�!�`�uv���x�υb��#�)W�gZOI��FXgY9S�u|��U�'~�$Ki�Y�y� M�z�T^R!*�/g 9��+W�uV�k��0��6*_m�It��ǒJ�w��l��UzN���u<����*
�{�dW/�zYk����,Ϥ�o�JM������'	.v���Gq������TbO��)�ue:�ޠi)�Ib����Eٞ;�I[Ɩ_��c�o������"���{YO�h�8�B��5W��^7
r��m���U0V�����(��KC�@l�n���}��Db7X��H�\6���1y�<uf�s����Ty'g�G�O�j�nŗۀ����
5��7��@��$/�&<�͘T$,�[A�`L�I�;�h%-p�c�-���%;���L"�7��p{9�q�r^ɫ̆��Y��)ǔ�B��NO�ͯ	|W�0��X�~��u��=�s �z?*���W7��7��β�;IО#/��t#ʖ�k��٘�%�m0�0�U
=6>aB���WϤ��*؀�ubk>����ZP�����ݝXƖL5���.+�z�(o	����Mjd�&6[!�R��Q�B�l��dv֎��;�������u�Nugׂ$D�.k����xp���#z��5��cbqQ��]��	��W�~,g���b+T�Q*u۪ź�}����y���
�_K�Z<��+�Ӣ�-�re�A��=)�xQ��]->A�Z��?���ۡ����X.+�!-<B���:}�*�Y�Mn)����D*a]S�I�#�QdG$���Nyt������/�n�#ؽ'���X|� ��u�*cq��ձ"��'��8�2��� �ڨ
geo��L�����9���� WGi�n:�����5v��(^|eqn��H�2%�.��*V�^H\�*���3�-+�p��FJx�P�FE�������HIҲ��%c��[�B�j���!���e4l1"�1޸x�CZ�(�G���g"%���B��a����"#��� $�����Yz��ve���#᳕L�����+�.�a�*���hM��c��d 1��.q�v�B?c�H��?�s�	(2 찦����BN��,� uL#�|ǃ���/�DK�.�,�h�ń�xw��|�`iu��7��X�
WPSq �t��Wa[^ֻ͆����S�<<H|i�'�5tK)���N�7���;=����J��8��;Z!?�uh��*��ρpK�J��ml��r�tL�Ȅd��dN������犻O��Pi��D1d�c~�
Dp��6�s�9��cz3��i��~������6�Fv��}]Zl��qb����˭!}o��G�Z{�rFj/��?�=ޓ�͓
��P�/�[}�d��&y-|�����hX��c����a���h*��v����҈q�L�??�XC)�1�C_U�!v�U >H��v�!�F� ��$�A��f�b�b���}yS�VGq�D"���P[�$(�Y�۾j�U��nFlab_�c�ԝ��?Y=К��p��=��R�7O��Whg{�X/�t��%`�C��{�8�L��r�]�F�C"'��Q\�ژT�x?�~�$Jq�L�3}�ؙT3�%r��2L�ŗ19CD����z�q�-�36�<��bm�r��	�IE���L�q5h�����߃^Z_�����w�u-�#T���`|�/�B�uO�Y߷�m����~�;J�@~���P�g|��\rbg��HZb�5��I�����x��U�z�U/0�g�*c�wg��&�eC����?Y��8a�y.F#Y		-3���rÉgέ�����==hyc���.�A�zV�.�6a�,C�&���@h�JG1^��!4���� ��<� �Ҕe��pv�_��eIc{�ڦp��jv`��Zܫ[�u�;FK��߬��U�44wMQ��2z>�������>���+�`Z>���ˠ����	�t'��tރ�ߐ���4,H+~F
�zf%����.���ng�=�%(0��<���.U�y��%m�^5�!rd�*����׌�?N6m��>���i�h|@e����̬|�q�S��J'���������0�N?�G�q��ʻ��냝 ~�8ސ3$�����UCis�C����^g��B��������@�Ut@ם-���b��?�Ð~n,қk�6�~>�|>;v�j3��3� yd��k��ώ F�'n��#l�(�oC����X�=�92�O�w�?�E�/;�)�fE�R��O��[�3Νåb��8�>h*�1��}S���@���W �����7/(V7.>�%�'�9�sE��K�2\�U�(�՝b8oU[�:&��{i����C.�C\�k$!]�I������|���d�G�U�&P:�Cs�S�W�4X��V+���WJ�%� 'B)�}B�@����S����_�P�GVwQ��F��
��%d[7���|�}~.գE�)zF�\��aa��9�������@n�z�/VE��̔<�zr�yope�6���������Ҝ+1�7Vx�E����fu�j,�E5���.W0󥐌bHb�6��m����mJ��}R�3�*z""{���%����*���LROa��hX����@�q7g?�Sò
���0
��B�e�5�u��=&��u_��v��R}G�!�$3O9���&bt_6����w����cc��ZEj�R%������$��
Ĩ���v��\��u�P[�R]�tk�Y5l�.��X�L�Nm�1��{���|yϴ�J��@J��tr(�%KuRب>��Z�0��{a�j�t�RI4�p���'�L�
|�G>�A���7=�����K�ɒW�����x�Su@��4�5N,��z���jo`�Ё)\����&y��88(t�2+���c�j�&;[���0[;<1�t6�*��/e�YYl�-Pw�����d9�n��f6��n�4�H3�$�CYV0��C�d�bg=��z�r`ፄ|ƭ��1#�����E#N��Ԣ\�?\��`k���JF�8�zY!A#��N=�iS���1L�3��D-��C���C7&�/�%��`x��j
�O���=�D�^1!h9��2/�P��bNV6
�����v��[�����[���{��O��B�U��b��f�؃$�3|��vַ�PR'i"�65ov|(���-��A��P!��UH��l���A@�����U ����R<}�1s�����g��o�V�s��{mE�kB��>�5B��OU��aM�	u�J�BRhi��c�4�
�;Ȅ�m?����'����U!3<'����YY<'o*Bj�� ��4#gˮ�u�}�$�v�\sZ�L!z,���6�]�=Z�4��Җ����5��R�eu��{�/�b �%˕��Ъm�z�@	�h��Z>�d������� }>��e�P���m/# F�%i�%��ޠV�X,*�|���mvO�L��l�J�	���d�p^��#�����:����埏6�Vq�]iB�|d:Nz4�L͔H	�c.y0ޡfw��:�}����C��A�U�]"����LP�5;�5�~>w�҇ �3�1^)�9�@.*�)�x$]������Tme)�{�vPSe�3idڰ�n!��Sd���P��/�o{��jҬ߃���a&���eB j�A��Nl�r���FEq��TW�O}U��������dy�龒�H����ŉ|�9jsǊ21��g�C��
,K"4p�Hc�4,�Z�� s�N��t�FB�F�?[&�d� M�#M�0C|�?&���D�M4X��\���@r����"����*g{�At��MjY����V��>~]�U�ټ1��wO"�e��(V�""Z�k���9g`
��pN�B4Hv�ި��$�U�3���W��~=>�b,���&���U�$�H��xC�3@��[	��j�r��^X�d�$�w��X�)�zd���B3]/�aeü�\�֖H4�7�KWؿ����g�����<0�1��w�v]��<Ø�0,�Vʺ��f���R�{���շ(ϥ��wb�*��-n�ϝ��Gߴ�z�6�<�Ӎ����9���̏�ׯ�3��ǥZa&T��ܷg�s2���#�!v#�c�`�ݩE�T_'�2(��`�����||y-��`��md�qJ�<E�� �ʰ�9Y/����t7�FÑ�ߘ;UC)�����/>f�B���	�I� ��֚n�`^�2�Ү�x�O_6m@���#�q*�ԭMT%�$�:eVY��6�0@k�"�6����Q�b�H�L�̠�J_3{�k�����@2��J7�J�/�W>�I�O�e�Z|cOi/{:D��_F;%
o�]L��z{*<��C�Ĩ>fo菭�7�ɨ��a6@0;jz�Ľ��Z7��g��N�bIXJ��FӆVVt��%��Fa��jA�GF�� ���O�E	�9��/���CFkG�ƕ7�Uu��E�=!�(�|�@8�ex����︐qK&-)̡#k�7�Db�;�0�4�r,�ׄ�'�Fc�]=���5E�ОV�(]~%z�m�����F��'9ɾ	����]W*����޼����}mf�2~����~�MPUYa� #����
F.��=+[����2Y�dB�%��he�ɞo+���1� N%����~����f{ ���}V��7�����mť]��m=
`�Lm�qÐ�4�����ӱ�M�:6��U'�/ڱ���`�;b�4� (D����F�F`s��GO,���V���U���p_�XTAf�������Ճh?S��I � K\>D6���	�`3��,eĝh�#���y��Z��*1��md�iW�Tz���_Ut���-����JG>�q��m�E�1z��@p+���V����E��z��m�Y*;r����刲�_�y�`Cg ���.4��I�-(lZ%��W&Q�rm�`�I\��+
��ۼ���}p�_!��C����&��]�H�|�h\�7.�fﺵ��`�n���9ʿ�jY�9\)��@y^j����<�oC�K�ܢ��1}ڤd���? �g�#��l�Fu�
�2s���1�w������yMtQ,���p	��TPtK:͘�5�I�!|�=�"]������7[k�֝���
�xv�|��Bמ��ӏ{*
n���_�AE�r���	u�߈����k��*e	?-�����%sΦ�mH	{��p?)��b��dx���+�+ۺ�-�H<��Z,j9*u��������P9�L��4�lx��C@=i�8�*3�*d�1σI�뙱GH���G^���nc��L�/�MZ�꙾6�'�7�9��/�!4��F"��6�=�mϺ\�xIǢW�2��NM��x��ߥ��x��&7�Sg�Ӻ�9~ـ�C0��X��1 ����`U��������,rzak ���o��6�b��qSh��a�b�TfߞR�.� �G��c�t�i�&~�yʝ�F�������3
)"
�O�@z�\,;�ńg�ܵ��]�������S"P~4�z	M�G�(��Seʝ,'*@>t�F���1A�읉].�x�[,kqWN�)�{��@j��
���:��4|���!l��Ľ���D���7l��/���k�l�p��lz�����
�֬�;�O����-�����H��J��*|Z}��C9giCH{(�ްj�rL�L��UY�P�����o4�L3��SsO���2�):��џה�l�sl9:�_��>��欳t��$&'��{�t��<w���k5IaP2��Ј=u���e[|a���Z���u��|�|w��癦��J���t��To��gn?��(Pぅ�K�ʿ�4��7k6��_D�ixZ�8IS#*dְ��?Υ%x� k�"��Q�vޮ ���P�������6���D�/�B�ۂ��Z� Cf��9J���s���A�i��w0���8?ҏ��B��/q���*,'龦�[�E(�n8� ��<�t#�W�7)�=-�&�
aQu
e):��τ5�|U��SZ��wD��t�c�	��S�>l��Q@���=�vɄ�6t��/1����r�����d{<b����CL?|B���Q����æԅ�'Y��0c����O�B��q�J���$W�0y+�_��05ه(�2�C�97"b	�f�5��RocI<�
1T���xP6��'�P0����eNW}���I+�n������N	�gf>�:�j1#���t�V�X�&x�*����x����4C��o-�<��-9_J�c�˭�`"1����B�O~���^R�UsF��c0��9�\�*No�hQ5k!�=y-?�7��/� �"KJ�Qi G���+Y�J��@�����9�}V;�A�f'W8g��HHg^{�wxm ��Q����Sh�Aߺȏu
��6�[V�ؖ_^�2���転�q�Ȥ�mZ�+��[6��d�>�R�õ����cV"�Gjx6�K�}Q��rٝ�D��B��"��X��{��SV�!��BZ��E��5}%�M�VWۇ��'�jH�p��q\GT�P��������y�`ߕ��j
����u%��2�xAܜiҽ��'�k���TG�����Z#�o{k����/���?�Ê`�n���wĩ��X����9���i��5�5e�c./�5ԍ��:�Pf�j��g\��<
�\�ʭ��m�}qL�Y�F�r���j�����M�����j�BO�U�a�2{8�g^]5�S�=0�C����r��JW�p1�w������zC��.��c�X��Ÿ�;�$V�-N̒��+���	ڜNr����K�Ǻ��H&*�8�2k�!�۶�XKK��gaO�����?D�����
p�nUFQ�]|@�+؝_4N�{<	n�4.�^�j�-%h~l◰��?�t�{G7���mt�����zp�ĝ�Ie�P	��>�&jr���;�!G� ��������Î!G������w����I`���A��x���r��|��+5�!w��u��v8L�s_�6�\����>�k������w~t_�Y����	M�bpƦ"����b��{��0E0K����Q+�j�f�E�*_���p��`na�Y�«���hF���M���`�r������sD�!>��n����F�a�<�m�[n<W��2b6j(ܟ��l��qGA���y�YA\|֩�_{UV�<J+	敟)$X��'%Z�~�\�Ya��-e��?P����fP�]�Devoe�*C��e����ׇ ���r�@AB����Q��ʚ�k����Meη,�`�����"����q�:Q�b���3��ױR�,s�p%u�}t{p!�FXQQ՝�Qx!�^��-yV��a�k�Jm��<u9�dNk�0v��W�2_�G�������m2���� 0n�+H7Ņ=;��B�ᓽov�8?A1~eRʃҋ���������y-��M3�Zm�*�u�Y�����5����[*����c$��U:�8`;۔�֤�a���(d2Ξ�1ΡZ��C`S�P�p\���[n/���\��H���¶IO�W��&Oט%��E!�b�z1Mڲ�M$������E��h%�kG�+LU�Hr&z��olcl�x������f���&�h��N�ږ^1��u���h�P�=S��3 h½�Bn�+ǈ '��ͣ�Kg�ٵ'���'c�Y4YF���~i$t�D�D5U�6Q�P���˜�u���D�f]K�������y|�	�:�̀: [�,���]��^��H�l3 0��}.���C��TV"�0;k�' z'�F��Lи��A;��o3�m�R�y��[�
�d��I�J$eX3�h6/Q�p�O��|�慤"��}��D�_�h�֩��Lv@�>��ڨ�3���2@�ee�ߦ"�pՈ���ޑΛ���c�i�j�#m�xֲWo�$�HX#{��O��Λ6�Ƃ�i2UP3��N�&����W��b(ZÙ�8��EJ�i�6m+�R�\�}f�@kۉ�>Z�����R��j䛱���n�<�7���,��*���k���n#RR��#Y��T1\�7N/�^Tϊ�^�n��6��^fU�y�P�J��y�/��mwGx�vdbU�5_qYl&jS�bzE �+�;Y7���l v�(Q��!��ȟ�1��=��@y�y��Y�g�t|-�W֤o���8�~֜`/)W��Kn�t���� -��
�g\�/uV���<�dn�tb��*p���{�Gu1����m���(�>��&��=��0]�����8�YUT���ϰu�Ln���+��AT��~�9 ���� �
�3b�E��e�Ȭ���^��]�ܻ�O��B�	��Z����q�<c9f,�Z�v@�GѿJ+�W)����#K��i�H�(�`=�י����I��z�/R�^V�<�Fc��>��t���$LM��$�6��)���H�<�z4p?�4b���Q>x���Z���,�G)�n(�o�:�N���L�v�'̌cfZO
n��ۏ1����PV`�*��q8H�w^�jEu'<[=+�p��1�K�s�Ϲr+�o<Xp��mr�d|�`��W`��N��Ļ/fp��[�
X���������ʗ=z�3ma8��*C�7U��(ل��1|Ԉ"�۽Y^m�z]��#�n�ZrF��� ��mZ~��oy `\xa��^j>+�[�@�����z�0r�{�ʓ (|��ơ��t���|4y��ϐ=�e��Vn�w�	�R9�BZ�k�O1$���9}����1��t����ȓ�V/���3RY����/�#ߢ�@�+�~����� _%;�C���-��0�1��HG��e��ٕ���s:z.�B�K��H�B����}�T�(wn*7@�ng�;e������^�S5�߷�H��E�Gՙ���>���t`$w�v�m�e��/I�$?��a�!�SJ��H"�?Z���U���⃾:�%{�^Fg��I\�,~-K�K�B��h`�`�d5�v�)"@��O����F���7�Jߎ����`���?~�;G��(G�ZT� �Y��s�?���z����&uZ\M��1����@�sSC��e�-s�!�qy�H�Vl6�ےbW���d7ūez�Z�Z{$���=��X�0Z��ҥ�pQ�U0d�p�V���������ح�� ;4����v����
K�?�D��'�����Y�{���;B�ui��Rn<QE��qhdDX<�lh�+����e�G�����2��n�(J�G��h���p�qC_d�m[oh��;��F��1�mj�IA:�����1�`0;�Q�:��"b��qv�E9ܨ��˼�)e�#X�]����<d�
<[��_�&,�W� �T�M�;��r�̊�e�q
!i%���ř�pP~�DX�-Y��pBO��S��

�N�<�q_74��W�����B��ԭ{�Ц�+���&�87�<68nl��4:����P4�D�=#��Ф����'P�Ҿ=/0)�^�8��\�[�֣~�k��2$7RVI�d��^��f zěc��&�8��յ��)�"���^>'w�"�\�Ɓf�N�FʽVH��P��Y�����Ҡ����?��TU�-)0�s��ѓ5Klqж������گ��1�2U<����N�� M� ���f�L�q+t��L�H\[N��4��_��~�o�,%C�ցZzvC�k~���yXr��.!:�X�������WM�`�VF���R�%9�g�<���Gp����<��\��e.�HnXs��F7O�M�؏тL�e���iYP�W�M�RI�c��-�
�1n����DR�2� ^~�?n�kNϛv��%l����@�n����D�\�=5��/o��߃=�|�s�-��6"^߱���m����2��woi�dH!$Jy�]N�z��3x�&����α�AGZ#�2]g"µn�(o��!&
�ϖ��ڧe�k`��Y����-'�k���$4\93���l}u
,]�}zM	�뎱h�*���X���7��i�X3|��+Δ�<s�c\Ѱ��}�|=��H񅓑-��:����aa`���sfm׿"�KvB�&W"����D,z �~��W���S����/�~3A R��� ���� �QV�\�$o=R ��Ne-�i�A�L|l�S�%�Կ=�9���PH,�qhU�̥��ɥ��~�g�4�<��${O���~OуlY3>��Z�dɿ%G��-���2�n�j��_/������oZ/_����:'ׯ��D>!�� �U���P�Kȩ��Y�Z�
���7}�[z"z!)Jf�Q}�?�)����Đ�a��W T����Q��i���c"���6�Y_=�B�(�e��k��"-��893g�a��7R��l�����pY���)<T�g{��Դ�	~�HG/qw*8���^�N}��Fb�����=}��}���C����b�ZjޜE���6��%���qI�$�\ԟ#;���u�A��Jh�;!�8H(-�4�b��q:�(B�\`��
��in�-18eZ���k��#���`���֮a�"�������1N��R}��Wa4�í��g�.����Q��d����?��9G��.̕� �h":R���.��&~9d��-�hz�v���L����L�rR�,��T����r�L�����}�v�w�iv}�{?���� �i����9�<P�0qD� W-�h� �O�׭B���Q���
�8T`�(�����.��J�n;��S����6�rd�-"�0%A}�a�a"ӝ�z�l�T}O�'?�#$�
�mp�2�",B�9����3�j5f߼->��&K��Nhr+���0%��^�X�f�l�%�1��[��4�a��g��;���~��~џmU�X�����a�S3�Q���J:q�t�~�`��D���L��|��=[_��ۈ��2sM��벂�A���PÚ<nS+���[�[ec3hm�#cxJ-��?Z�|B� �*��߽�z���n��9n��.Қ�O��r��V?���V��_-޸eu���f&����,�*xKeZQ639j$֊J'�ݯA�u��ϕI����~��9����L9M~��]��Y}��4S��:��n��B����N��	|����Y�nH#��ҳ�x�֞߼2?�I�f�<�$��͜�(����h�ط��le��n�n�Z`�r
�+R���(W��gm���B��`����dٝd�9�b�%�G�Tϵ���A�P��F?$H�f.������������JY��Ow
VH�8(i7X�j���X��lQ^�����WJ��oMC�Þ�GqK0h�X(�{�5��7������[�M�,���^B)��<�r� ��z�4��b&"���'8[��X�>�$w���I.��7�-w<���!�Πla��91P����
�|B�8��t?zz03/�s7��ni�0ޜ�Xg�켛	ӇL_��J�M�������ӄ_�+��e����L�l����XI�ǈ�U�Y
�n�����}YD<�<;�N�=}��Ĺ�����a��N�8{P2�S���D��^/SSO���� �#l�e(&L���U%�Q��_kp*D����(`�7*�[�Q֔0�i'�QY1j�v3��I�Jp����T��]��M�h�h���"&-���BT��)��ϙm*��@�I܀O��F9˃�ߢ<I��a �x�	q�fH������ÕVwE�x)/�\v�Y%�����)�ޅ�~��taC�Ȥ�D+2&�n$���B���s��\��N��%��{Y��L�?��Ja����:�OG��w���r��+Y�b�МLc��Ws�iC���ӌQr&���m�,�P'(Y���8�=r!���DP�Z��&]�H�q�Y};����a��jJ��`Eh�SQZ:�)EM�v�L�5�l�y��2&�߿���є�%DR�RҞ�J���XZ�to�l��� g�4 7z�.� �q(b�yL�����Wַ��(pQ��85�`s��ꁞ@;^�����(���~�������[�\ʰ7mYS�Ԫ�u6H����F�0b��ɱ��ǝ�қ��~a���L���;����<�l`M��/�G���D-�+E&O{y����f�3>��pga|!@7��]?�;�,h����7�l���#�G\�`��q~��td䦝M��h� ����9�n\������=�¢hl�ӕ����Q��q��G�%^��z|O�ٍ��~/��n�[;%�z�N:
K�x�:��9<��Y�Z�X[(�֠9�����?>��?9hB/����$�J��:�ƞI�(J�b����X�'�!�k:�L>�)��bϝ�ma���	
�Ԧ������aI���Dw��Yé��t[U���>,Ϳm�E�k�F+͍�޸nɊ�q/�MN}O�s���9C_���5�1N\�N1b�aT�D�ae��}*w���ા�N{J*�8����`�V�J���]�Y)fX�1� V�����Q�q��Ҹ2>�|�R�i҅l�D�#�~׼�=���Ϥ+=�Vu�va��m�闸5���1���W�c�w���E����w[#�� q:]��)�Dot���J8�׹p�N��H1�O��?�"ܑ��	�}�/+�Fd��c�t�k�q��5��W*�a��ʼ�t�����F|��7H�0���Y@�&Rv��b�g[�KlYp3��ޢ�A�U6���Wq��-]�pcs���"p�3<��y�9k�X�q+�ٙ̉"o�<m��3̘�4U�X�CК�@4߸>��9�f�<���V_�A#I�â���
��R�gIc��HX�ˠ��w���J��{a�����1�����d��-�<��	��.Z���+�ˡ_$��9
0������3�D�fH�S�Y&ⱥ��L�:ٺ~O��so���п,uOo���I6N[M1R�Sx��94��qۃ�E�SN��Y��z��Ñ8Չ!��qگ��y�Q<����+	�	#��?"5�̟�<��D@�JH;-���==O�em����tP	�8��@xϙϨ��k�����j��[!G9�o�����MD��a�V��]���<ZI�@zz$���NTE���i��"�H$�uFD��W'#��w��ۢ���$3�r� ��U��誁E�#���.�tɇ�OVD����|�Ѭh��m}��a0�����en
�״'�nK�ud���zRX�x�+��_:W�q�5@��d~ +ʜ�Ou}����1�چ��( Q@�f�R�P9�篊p�ĦkѼ�	}֏�� u���j����'zW���_0����o�c���7N���(nCgp�R�k���Ւ�Q����g��S,�$����ߖ̵D�����_�^���s�y����0�"��ާ\��ss%X�Dz��qX�$Y��E:�*7?��8��<4S�;j��T�@>�"B�5�L��ϴ}g_b������n�X�2��}?���b�~9"��!zH����P���}�H��h���a�����ۙ�/}5��jW���<_2��V a{DlX�����&�]{4��м�B�u=:u��;n�8�
�;�VS��{�^�U8�P�pJ�B�����|s����Uc%��
����e�#}+�{7�bP�)4�R�������y���	\{g����Y��F ���G�.�l=�%������;w�ރ��`{�{NH��ó���H/NT�̤Y��:(�Ap�;!��1�Cȥ%��f�
�P���]��:�+�IZ��[�bsT�s���|�y3��!���c7/��_��U%֐(��8����2"ݺ���Ӿ������o�����i�ٲ+5�K�Ԁ{�V@ܽV���4� �.}��}�:8�Ҍ����ɿϊH�E���)9=�Z����*H�Y�qWJ(��� ���1�0"���ǯ���WC&���a2�������u o(Տ?@�!�%�}���ȵ�	��Y��?U����.uz��Me��r'�+��o��٠��RBQDvv��{[�.2�����pן����F��jFt?�.�̔W�h�mL���NeJ=M�	��1�J>��U,�m��6�����̠��ꑲ�11N�[U��ȅ�ƥR���=���B��=�/7�ズ�O<(;k�Cġ�)��@�*%2���~�k%�1�z�>h���LB��.����d��X��	,����h�"y2T���p��������+np�O������rc��6�қ�s�Vn���Mb����m�&}��^M�١� �վ<�0]�o
N�ʄ�>��M"+��K9}�rSX�%8�\�Wգ�|b�O�̹�^��jBG�d�?g����������,�OsT�X�J yw���[I����( �#G����xd!�F�f��N���`�\�s_�u%v,�!��Ĥ:�����X�����Ɏ�-���0x ��\x���gM����yY�e��C��a��{a�C�3��ez°��1�jxb_A��Qb�ۯ�7j՛ˌDިY�\�|�a4��W��&�/BK�۲�Y|p8��n`%hY-��T�����m@�鱠�`��y<�|5D��)=-���8�V��6�֩ج�������)��F6{�l}�|`�)v���=�������`[�@�D�Lŕ�5r��ʦW��{)3Y4.�8鮣�3nSYf;��>�w�xf<[&X>)�ñ�R�G~7�z�}�k&��`V�%�M��0���>��r�@O����\����IxUOѐ���|�W���� �&�b�3��:�Rm���7�k�����3�� />�"Q(����~0L7_��T���!��f�c�B+t��*]"%D�bo�оs$Q7�?�*��b	��ͩD>4Rv�����J���	Q�J��2�j��U]�D$�����RU��Re7��Ӑ�w�N�#������Eyo*�'G/�C������V��)�oߑ:��#Y�@ۊ/������9�F����D�|�r���2�����niV�g��Q�_����ub����}�v�d�J�o|�2���̤�l�Q4t����ޤ�E�
���dc��^��Y�����آi�CK~&��i�[JL�V��8 �ˉm
��0d��nٚ|5��Imv��n��5���ڼ�L�Ԇ���@���ad2����o��:I=�ڬ'�B���X�>ӣ�������ɆJSs�,L71<��K�k��*,��hjK>�
�i�x�����+r90��VP}6�y"�ls��8p��O;wdU�9.����T����=;�b�S�6�aF'��lʰ]��ܡ1�hJz��N�id�5y�����m_���B��(%��!g�:�6�'����vMT|���#��ҧ!��\���{�� ��]S�'�{+.t����^��k�a������^���3�nB��_уk�R�-w�`�.�Q��ɯ+�M���LW�^�/c�iT�� ��y#L��#58S/����uAH	��J^۽��s��[m������z��C8@5���c6;3���,�U�y�_U��ؗҼ�����g����;��D�i��U�V�7�kc�|�ӻ��.�&��O�K��zRݫ��!�u�.�K��uD����A����#�?�Z�b͌�\��̨z{>ߵ~O�Q&(�S���׹Z,`2�賈���J�4�/F�r!M�;�ѻ�
e��:�0�bEmFJA�G@�#%�ڂBl�c0xڕj<or��V0�K_l)����)/TG����:鉁:�T��/^_�;}p�[�ˢw���=\�QKy�D�]Mג����-:�!��U���	]
�]��%�p��c���`���=��_��e��6�c�Ƕ,���OJ�r�Ԁ�l@�i9�����]��BI�K�E���)s�B"/��I��|J�>�ˇ�Ͳ�We���3�Jr�~!�Q�j�u]]��Yy�R ���n�-�1�dk�m���'t﷔!�S��>E��I�Sn�ƹ�S�1�[�@��\ �6rN!�1��9�Q�ͺ��=C�o������U&󐉣/PM��vӖts�f�U��e�W�/�~�d�G`A��_b���{5�Y
�ah-������ qBsLA�NApL���$
����;8�3���J9�$\����7Ez��������k\�����#�>�߅�Q��,��V�hG�f�:O���N|�S&i��?����X�d�Iw�\����NVO���K>��|�<F���R�~e����)�5𭺵ּ�HmB����1��H>�H�n�;B���2��&�x	��v2�vS\���c$O������)������5'8�w�����:L�v�>I	���ᐄ�V��쟰.�ʇ�͠u�m�YK�����:,���ܻ�i��4I�����\7�s���Dp���t����Ti� O���VJ�_ ��ac�Bkw�����0H��h�	��Ӫ���!�20���������9J�1��KaB.i�\1/�Od0�4�>�pY��9�d���IT��
�p���ӫ#�~���\RP�����,�O`fQS����E
�z'��Q��pww�W�9Y.�Ru�%Hބm� ��Ŷ]��BT�"��Z�_ ��2�=t��]M���#�o^,��w�xf�Qz&�6� �4vD��p88*W^VQ�쪎Y�0�y@aO����4���ꄾ��9������R�c�腒�L���B��R�4��J�+��Ӂ$c��$�����c_�$�x.��JaA8&||�������R�v�>�;���jP�^Q+kݖp�}uܟ�=r˷�L���E��6�y�X�J��}�|�fL��"�ŝ�İp?��j�G`ː(�Zc�E�W�Bp���<���T'C��-��1�"�Z���Ä�r i �z�T��6���S�97���Te��&�]
ͩ��J/=!����������MHϻ�D�h@"�d-<�o�F�V�+��zʁ����Պ�l�����i��&��Z���;�eԍu�KH:�@�+I�PG�����B�z �V�F��*�_���0J���� �1 {^�"�/�q��)���oV��T-�F!S �م×{�ЯPD*�9D:�n�}�{�ӟ.�M�jz�\A� 
�g1�e �ǖ����^����фn�7����v���F[��N���n�3é֢� y���c�b54Ȑ۫4�I���|� Q4���������e25��S
׳+��V<CYZ�;:?S'�L^�����B�9`i(���d�`JG7\��[�MWI(y��D���DFj�ͽ;�,ZM���.3\Nx���I����W��D&	�H4s�����8�)xүK'�6T$�~�2�a�K�Θē�����ۡ�P��o[��ki$Ή�����I�ۘD�l�1�͠o��`@B"a\�Hܛ�VpM�[����@_�����
@LΥ�T���7����7�3I�D�H��'��1�o^j�������'K���yh<��y�D���S��%��˱*ߤ�i���2X�Z˼��'p�J�[yVj!P�V1��OR4;��Պ6��TR�g������x�h�W����)<����8�r��(��O8n;�"H�DŹ��Йنt;M73����L$��kt�!��{���fr�L��CZ4�\�d�:�A��a�����Sݰ��4Ej�b_��	�V�6�V�8}�i:SY�O�ӊ~B�p���{B��T�ظF	��Ĕ֐�W������}�$)�g֦�9T9�NeP�^+�d���洗ꅢ"�4�c��([��)MY�+�H�,GuE�l=��i��[���8>�*�R��;Kyv�F�d���L�� �;b�"�dy��y��f�ԝ�8u4/?��a��̊.���&�6��)�m����'	x�[���d/|jJ����NP�'��Ǆ�xa����	g5xW)x}�X��1QKS|�nA��?|B.W��M�|3�L�������4z��$�X��aў�M��ӗ�r��wQd�x�w87�h�U�HA�m`4�;���=`A.y_≉�&�9	sp1� s���Ӣt��p{P�"p�����E��lz�ȼ���@��u��E�JH���/LR�^	ݽN#D[�yZ��-���{��)�m�x��L�	�s�捘}�.�����~�1�!߀�-���������E<Z��,/E'�`)ǎ{�p��r*��VСZ��q~t��`W�2﮳r�wB��c��z�»���O�2]�j� /�R�x:��\iLD���5 3�Hȣ������A9�b��:�f�6��U�PlF��7��W��-ӊ��A�D���D�S8(O,#���Q{=\(��[�e�ͽb�/ ���`�w�10�xj�9�R��q���swb0���=���ڄ{���)������O|vc�j$dd�E��|ّ`3$��s@�c�iK	�R��i�ݚ�>Bկqp��?r�0���
З�|!��f�Z9��_Lf��p.@�B�g����"=HJ�?�1�t�: �ۜҽ(#v�ƺ�b�l�����n�m�϶���?y��"B���_sѽT�/�mM_���CɷJh�=y��#�&r_r����-�Z钁-#�������j��Y]A4�"�r#���*��d� 7�c�)V�`V-�����n��ȮBk�ֈ�N��^� ��U�|I��@�P�EM�19�  $��P��S,�%�{�S��ۑ�Tc��dҐ&l�æ�*��Y�Z.{�G�j��z؊Ђ��슧����,�]�/�c1�ą+��#��wŁ|R4�D��nɘ�n��0�]�
�&(0���k7�� ��C=�f�4��_��I�{��S 4}`ʜR�g�m�uT9}r?lLA���u���7L?����1=�����y�l���Zse@��>s����ݰ)G9]y���uK�
K$G.}�'��#/z�]O�l�U����y�5�6{}R�{Ó�}����Q1���vA~/�qxtr]B8�Ɛ�?�y+n���������K���N4�Edh%����sib��c�L��i1��y�R�(�A ����=����Z{�/��;gRA�;@֊C�����5�>=0�-�vִJ�����d���ۦ�]�b	E�,���8��c���H������Bt�\��.-��F+�r�Y������|��kg���E��xb�q����[��Eg��;�a��`�&Q�Ng4� wbS��@ϓ��-��c��*�O&/��_�Ȩo	)W�,0��?�ͪXC��̳r��a�;�0��,f��*��ǅ��u���ϻ�ZI*?��R(��>��o"��xV���������ۯmf��\[1�M��`�;�T�B��]�l>@��^GQx�������G�}�DrL�G��N���Ɲ�Ra[&�z,���0���q5�Jޮ'��>�:�>��1�R&�b#�f��,7�3SVp�/�D� ��4���|k��P��qAm}��Њ������>����m������Y*}�)@�)��^i�����9��H�q������ RF�S!a!�g0��ٷ^�t�!��=�zmPz]Lj%���e�<z�ʴ�"��'�z)�ӯP)[P@���o���7n��&�������f5��	����Ve���A_3��9��\��i!yw�|>c�����#��ű؜�5��W!6��]((�H���v�J�I�4�b�w]�L���ÏDeP�5j��^0�^�}�r0�8]��덬����V���d\w�NA�L���j� ����[��Bw`�V��t?JN��#+�c?K^��х���Кj!n_�:~v�\H9��S�=���t��"��� j�����Ԗ��.u��r���5�|�������n&w\�rN��L=��Nq�u�
?'���g��ӷl�F�����)��B���0�Uܸ���N�kSl�ͨ��Fx�n��RW�]"��i�ڠ������o��U���,u�qZ=c��/8�[�+��G;�PM����N�Ř�H��
���|D @x��=�=�븨ԩE��4Wc��;)\�l�����ڐ�*�"�n��z�p�d�2 �w�S��͓��Ѣ(j�AX"�i`�b)
.z纉�;"O��ֲ�,fC	�m��D��{��$	��4}���]���AУDh�L�'K� �ǲ�*N����,;���jSp��~���"�"�jx5&~۴3��S���k£u��23����$p�%�1���~e+� �AG�UGl�.��i`n��񲮥�P^u��a��u��Ri6Z0s�/+p�z�����r%�?*8��0�$BB�:�Q0�:�/	��]����K��;	m��@��`���zO�'}'(�	r0{I���r�ț2��S��m�W�PET[�Ks%_[����t�!]��oň�áR�>�o�_ȤB73!���)�Ыtx*��R_7���(�w�n-B|�-,t)>)�(r����K�eNsw�����3���Z7��NF w��4�(���[�P撉}��
a���]�sYKZ�I��-�$�%n�x!���h���S$�L8A�%���!��W����{�����L�jK���k�`���l��t����OV�]ɛ3Z �d�vg�Tkɼ\�ә���%��g�'����Z��t�,�b�1T&J> F����E�O��J;�4Z��A��d̓��*c&g��oӅ���攡El��n/����;r?��S�I���9��V�:!kexv2/|�K��qFְ����6����G�y�#=�[T�g���KM��V9��S	����M�$H�U�m��b/�0O2|������_�RS6b~�M�N|sMRK5���+��!���KN\xBK�E4W���1�N�'�e�$�~�J{�8��{���h�b�T��$)@Ɣ$RP�5�D	"����i7,#g�D�0��V!Z���K���Tn
V�1EFUK-.i=�6l܁�(ry�V(E��G�|]�@���["��t#�݄��� )���qGvA��(�Ǻ
e�I²�,�1�)z����љ�P=K���7�~��"���J�=+�.����VZ�/�]3�L�}��^����NLH�E��C���%�J!�cY��\F�Nԟ��s��n`�� V�<�?p�MM�=:����K:�<.�Q�g�&&��c\s����O3l?��M�jEoB�@}���>�	��ߠ�� /��HI斧��zH�$@�ߥ!�h��j!C�������S���m[�[�sĭ1��0�9Wa(�,`�F+1N��2�-P�F��� uC�ڡ�""�3���
�ه�[w�+08Y���������lI�)Ri4�/�G@yx2�)����M�J��d�\U�6�||�t��m��?�P�`1���,�lC���
��|��|�z�"#��)	zf^�!6�ft,O�2���4���ՎR�ә�+0f(���-��-l3Vkot,;��P�=ۊ	���w!�b:T��@�=��5
�O��è�u����RU�9��e�fGz~�k𸚚=�����
쫪�����O���}@��Y�1r3 � 6.�����h1���L�x,O v.I$z�R�@ɞ����CJ��	�9�r�Ik*q0��2�w�˫I��<<̪z��L��B�mL[J���)TI�D-���0�&Y@�g���@'�-��nN�����KT8��.Ϳ��pʜuwjSF�?���\5҆N؉�J�PO��Kg)�J"EMn ���W�O�=� �G�4 �an�6�"&��:^�3�E9!6�%�-��GWAo
�#҆�����h�V	|W��SfNL>P��8�� �����pq�-��pc�W;&�)��{��{\��6��YୟM��M��;��h�Y�p��p��8֔=-6{����u���l�W����S���x�@G�!~��&?�f��_)�ۡ� ��LkI�*I�	���}8-Šx/I�[�-��\X1�������.~Z���u��Oz�a�@�����(� �^�<�d�?�F+Lc1B���3W��dz�Ms��N��H��H�b��e�uc��q*���>�hǇ����/��_�c�du��|�P����Up��qV3075$16;o?�L`�
\�K��t�HA�Γ\=L�魉��[�\���q�Z����8c��K�\z�ylI�
�MlH�և��c�%�FT/���G=�:ڏ�CeW�CO�B� ~h(oϭ/�^m�!T���?]~Ү������BoA\y����,Z �h1^�����OkZ�`�|��k�[�psr:=�c��]�G%�
��}<a]�D�퐈��A1��8^�X�گ�)��~��n@$�3hw����?��n�H��Baf�bm:B3�N��A�o�����.���P�m}s�"��oBJP�[�UZ�x�@ҡ���ts-�ٷ�g0���]R�Dz��:��Y�I��e޾�z�����׽چO
�{��7}�2?�##��'���MBw6�tU���'�
R(r�ł#q�Zz�q�g劵J[�ӹ�Oz���3�v��u��C���O����u�7u�d���.��`>�&��sv�]r����7!�)���s^N.�T�`���O]3��Zdaf5]x�o��W����9��=9���q	J��7DI��W��g��D����d�@^��/�B�V
�9O����C:�η{���/>"���mP�"����h��3o������{���<�f/�K#�`c�s_��"�䍄�jv��s��-�M� �JW������@^�ck�zu��Lë�WQ�� ���7J���V�G�K��[mo����0j�7b\|�$��3x���q��n�,���sr�:��r&��W��Y;1�6 ��P<���e����eZ��T�O,�q�����L|��M�G Y�dj����wӎ`A-���-C�8�%��4`��j���	RP#�tNM�hm~��ձ�a�䲢Bȴ?���ܖ�o����{��`���؛��d�^�+��$����z������
�y#��4E[���=���bDى�N��fˤ��񾘷����qw~�*��hFZkUQ��H��7�M�!���YU�Ã�:�a_G��6˺ν~
�Ֆ%wm2m�����Uoܠ��<�������&_ׂ���Ԛ��)�o9@�gNYd��*+�"�g#�y0z1�p������N��7L܃�#|����rQ�1���݈�
����o�É�����Nd�n��/_h��T_�H5a�WB�W[�b�o&�f�}\V�  ��"���c~�4�`��"�X���2���V�Ƶ�EЫ�h��et��t?5^�
�w
.�� 7zK�쐧7��sa[N��>��k� E�j�+�j. �@+�T�n�daYre�)C���������~y:��
;k��j�ZՆ�Sk1�l��� @'����9�C��ZJ�8�,��h��0�qJ��'�AY��h��q<3L_�S��*���Nv����N� ��h�͈��&��%uv̖s�E�V���1��vy!�,�=�tÊfN�:��"�n�TA����d\[��'�o�\"��Y�z	)f��TDu<j.�qל�Y�~�]=�,�&�A7��}����Lh�8{�`�7������b�j�1����ŏ����H�1�}�_F�0�a^��/[�|���R�����P��/F,$ ��̭gv�I�t�/��[J3�
- �4}���<���&U��
�aRxa-Ā	��6`Yz<�`��8�A��f	3���r��2�x�o{��34���~�A����ߵ*SM�@#k�_z��.�������z����׉A��D{�J�� ��R~-����?����]�������ؒ?�_-���G;�x3�zuD͒q��$������V�cYD�;��6RwI ������-@����,j+|h܊N`g)Ɗ� ����j8щ�&�A����&���~���#��$73�BC�~gƘ��ܐ�V������$�٠�9!(FF�f.x�y���X*2</��Ј���̆���=5�\5�B�"�ʡ
t��Z-�C�1���|��Sk�[C��Z)h��Š�z ��{���vg�>�]r��x]�R�F��)�\�*HH"�ƦF��Z*���;�[ii�틀
xpn���2�1Z�x횬u7�H*��7��k��t
��#���9�51����S/蔅k�<������Q��'x���_����:%㫊A� �� �G����&䂩���{֙9�"J��3	I�n}d_��^9�������a4d��unA��sQ�'o�O��`}�EW�ӂ~��6�}����N�3W�SUM�;q�`NHC>`��y���j��Tv��6J\%�o@S]54Ь"�u�*0}�!37N�a䤞��U�i$�h�`�!$xzB��/������;ҷ�����l���l�"���e�h�NUrS�Wm�%mT��� 5���z}�����RP���`���b�ȃ�"��|!#K'rf�&�U��ó��MF*��w�n�K��֘U�9'�y�Ԕ��o�~���k�\"�;�K��F�ȗ��]OHnf#�S�i�����z�*M{T֒�*u{���R
�F2�z��i�� S����a��2,�
����f���7�6�ѯpD����jݢ�Jݹ1�b�9�|����8���?DN 3�Տ>&��=N��[=w�R�@;[�6aд��kt۠��yt��GHK��P�_Z�����xt\�v��r����������C=�&�ד�H[Y��̉�K� 3D!���c�a	BF�?m�iǫ�=��^�[�>ײ��� mCb�8k�+8<�j�-�����iS>nd� ��2�O�Wo�D}B���1�.�K7�ǯ8OY#��Y������2mD�z�c�ב��6��l������t��'<ne˥�s�Zv2�bu�m��w�1�iGOO까sD�Y��P.�zY��y���Q�����鍢����JP!/�\��ZϮ��^}�#�%��p�͓�f�ނ^����-�z�}����t��ar�lL���`���ƥ�^�~B�q�����5K�)�\�[\�a��-ե�ΎK���/^�����<��&g�sq����d���4Ց�!���}���!�?��[OB�{VRܤ�B���0T�0�BpC��%�oȟO�?GR��K��=Ҫ��gZx$`������|� �����S5H���U�NK�z]y�J��`f��-��r�U���+2��4��Z?p��}$�|�As���ιL4)�l+ {踔׳�+YuD[wn��M[��	���Q�خ2xoĽ:0��Y�W��,�J��#T�����r37���`���x�2��I[�'�+�tꫛ:"B4�X�^��꧝.yP�X�\v�Ϻ�i����	��DL���d�����V�YC!2`Ca�%�=i�<#��ʻ��
8������2 �!�x�{~zo���.`�ª���k�i0Ews��;^��G+/�	�P����*f?��J��m����<~~-�C��O��7�Vj�60�E"�;b�e,=��#�m�lo��e�ܨ��wq�S0)4T�_J+��.�\V�ƥ�x`~-��o�nl�v��_�/eߦ*��.�}����C.�\���\X��X?��`�����z@��k%]�@̥@m&���C�O�0Qh ���T$>l�cK8��
��	J�;��>sk3����jX�'��Lo��)3�{��U.w�X��0Cg6��$��C �=F'�>	�~�?�6m	º�I�<��*7~�]��p/,�&����Ѿؑi{���0)�������&��t�caG#U�TT���i�E2���}�P��c���#{#�Ζ�u_�ʹ�5r�/ݨ��ܕ��Ȭ��C����>u�B��H�J��~�=<o3#�+��'��k�j�xze"]ke�=q�O;H���[�uZ$������T��E��l#\�so���T
�p��@@P����@��L�	&pM��aB�F�0 �k��kl&o�u�����Z|�r� �*�ɸ�0)�_�)/��ԣ�������&h[fd�Ì*?�g�N�b����]Ǆ���o�b֘5ZB��<��\��RS�t�p��:TeN��%��q�9b^$�}���G�k�$Ov��y8v+߭j��/�mN�o6�����(=*�s���Ϯl�v���!(�Ԫ}%6`���������c���q���c���]�R��e����ߓ/�%�:�}~��Y��Ա��8�V���m��
�Lȍv?�[�<ϻ���v&Lh��>�p������G�-E�9��[Ca�6e�������ы�����)#,���5敧;g�JzL��RǶ\	s����kC��
�O�����{\����Q�	��(l���c\�_C��춹)&F\�OJ�Oș��֐fB��[�gc��h5y���XjW�r��km
�u븾��n��y�pK��Z+�\��)&���y/۷?��ڷ�e˕ Q}t;�G���v�d�1E>��R�Z`Lakp�܀`�j8��#z��ɜ-{����y�A��2 F���i�HȀ�c����H��ys*J���r��q�$%��ڪ�^jh��lkc��%��͚���&Dx6OQ�D�6�fH?���ʩ��t
�j�?�F��]��͓��
��v��~� ���x����=E�����	hݲ���m�H;��T,���Ov�6���?�	��i�m��bG	���[�x^��)a���I^^��+��3ˡҞ���U,�m^������u��,H�C:�S5��M��jR�g%�T��sf��E<o�M	a����7cc�'K�f6KӢ�W�^
E�&;^��C���Z����k˙��O��S	�z0�}Hx�r��g�N���-�S��ٰ_���-��E��J�a�4�h`�o�|Yz��ȋ�IJT���/���h:��]���cBP{�ar�+?����/������el�Ѩ�\��d\�U<�H�מ��d��y{�F���~d��w��I���:a�dp�m񯁝�Ԧ��z��`�b�X̎�҄����*����8��S�9�F�h�k��	��8��Q�8[p���P����V�G�<�e�xj3$}���;QRט�Ȓ��Jv�q�y�^+��:@q����$}ޗ}�^�xx�s`ٶI�H�T���Ag�W" �H�H���� j6-�^�{UZ������7�>�/�f:��^�Uj�;BR�Wr�͉��u1^����;���;&ɯ��,g8���ϒ���ќ�����d�v��l��r
�͏r=�8�wWb5�S��H�\��H/�K�A+n����]DR�
����)mv}�ʛ�!��`��6�����.Cb)��c�� k@����5�C�[�����8�T�ۏ�q&�	cz��c���r= ��<����yES���>�XD��%�� v�u���L���2��-���'~�=[�;�(�8�8c�����Q�<f��'QY�c���Ʀ�>'���X�t�%�	<:���|�.}���ך�ﲩ�[��`�<��Ƃ��R	�!�m5�d%AX�XVHxf��sK��"gσū���Rx��G�X=�d�j�%�\����X� �P�fc�$�.���a���F���G�h]䜥������N�xj��d�zP��7�-�K�1%޳/���q��Ň	7�Aj'��߃�0 I�}(Q����&�Yf9 �S�!�J�D2 0*�8�[�J�yk�6e���@�i�4�I~�����g�㈮�y��L1�l6!��a���F)�43��S'>�/L����^�&�1�s��U�ptp�&j��!F��k�O�f9z��D���g����F&MX��gI$�\H0QD<D�ؘF���wV�͉/&#��ӝ�	�!��֒/�RC�{{η㛆�9;'3JA	��5�1��b��s�Z�:5	0���6��>��<����Cb#�g����6�.��O�@7x��ח3��k;��nD0�x.����O�(����� giN��"��t��m}�F��د6��Ot�+��d������Y�w��i:~s��",�*,^o������Ċs[3�K�9��j���{���˯������Բ� �Ȳ�w���|��u�)��!YE�#;��};�k�D��\�9?=#�>J�ޯ.n��D��<��GoU�G��<��p�
	�A�������|P+ �y���Jk�k��*;1��06.�S��ʕe��=Û�C�%.sW�W��M
���bE�oz�NJ�3�I]��z7>~d�\Q,����d���#oT�t�hV8� wn�Z ����^�r
�cZ˺3QG2Jr�pmo�&�I�k�܉_�sGRz��bX�N4�O�sw��r��6�rX���찍�$K��cr�~}�G�[�������>�0B~\L�)������4�����uE���﹎���Ym�	 ��j	��ʪ��'lw�U;+���S/A���S��Ȭn/Y(c�?��__���{��2"/�����4��V�N�	<����_�H�$c�����?��y0����=�Z䐤��%���wm���:{�Y��rj�4N��bRJ#R}��Y�H ŵ�R��7dˎ��o�J`��!R�2�a��&U�9�ک��:�1.����^�:M�8�NH��0G| �ɱ�ºIO1i�X�K�%�ݬ�ꂗ(�����=��������z��J�qdТ��}�-��1|���M}hW�nh&oc�0os9r�p8�<7��~]��k�����5NB��&K���/b�H3���/U��^{�$|Z���בI=�`$�p`{VU�W�XIB�X��}�ʾ��uw����J��ޤ/d~��h��s����������#��&�����Ek����\�-�=P��l�م
å�mϸ|��Й���]'����7��C�=��m�Q  ���ҫ���OƖ��"u��ʖ(-�l����c�q��ƨ�mhRL���%M@��Kq��- �]QQ��q?����#YZ�V�����i�qWTm�o;��8#/A�
I�̻�7���t�NY�c���Ē
��K\;Q��d^�i�G@AG���e���wOt/�$�j�������&��]�7�-�6������ke�p��7{�T���eVqcNw�v��l�u ��#7�#�o�P�؟��!Vg��D�-��J�`KJg��z�N�O(Q�V�@uW)��hNBG�|�-?����:UI����Z�*5�<	��h-�U-rq;-D.\�4��M\��H�Z~���O��㎤�٣���Zz<���RN��沦k���õ���9���>'%<%e{��b/Q��L���W I9�MS��X�w�"��/Y9t�B�g�lUF9T+�c�����?fZ�2X�7��@Tٻqw�����)続��З�r�#Q|���R�Mf�2��Ȟ���U�&S��K��[R�h�:��v�ho��[��fPq���	�U�!���L-���������йIuG�z�Fz����Ȩ,x���ч�n[�����CN݄�߯+%|�M4�R`��֍�8>�vh%�j��#ڥ���j�pǇ$%&��>%��ˣ�L%�j�42A�)|/���D��CE:۪C�VY�Ɣ��0+�����	���B�1�5<c�Љ��QO�5�F_�~1w�&�@6�=ַS%��6�qc�g�=���dt��A|�v,n*�ݼ<���U��D��������εЁc`p�a��2ٙ���������=���~��LJ��T�L�1�J
d�OR���ۊc�p�py��ps������[)1��;AP�k�T��:���yN�I������ĨJ�V�2)�,���o�����X�<�g�hNj�H()>���cLw4oK���t}G �����6.1�(g*�DQ����R&���`'Z � m�Ӣ���&���ɳ�7������}��� ߝ�=��
H����BI'}jCtmcN����x���y�Vj'Ԣ��FX����Dڢ��~���j�'>N=�[~t>\�r}��d��N�D1sn������{�Ӡ��K�Sj۩�痃�ڰ�}b���ҫ)ǵ�/�W ]���~��.���K�1C�7�=��������v�B�%�0���9Cm���Yh`D�\W�Ag8��HA½d+������Jc}��Ტ+�	�RǈS �kI^�
��@�=��j2�By޶A,.��Wa\���,F�\���h�Ig^f4*�"B��3��ů��G`�R���8��7��Z\�''���'�G?(�:Y���d�z%8�0N��D��M"udQ��]�6�j� ��L�R�%9��7��d'���Y��o�"MT�H��K�`O�A �˗�d�E��`�Е2�琘)��������`�O�«`Igcr���58�CF�Ù��9~�(�X�1���7HN���S\���q��႒)�b@���(Y:j�+6Kc	������$j�+��m�;��7\�^��Lx���|V�/���CáI�Q%C�iu�p�TjܩŲD�_+$%��c��]�h�0�Y����r�du�� o�Z�Y /̃Y�s����?���]wCų]��w����s�M���tk�鉅ld}/S)�׏,��L5 �afDb�ء���|�p��&�5}=����9�`�)���o�0���h�L�<Rd�
!�X>����%�a��,V��k~���x�w�Dy�K�j����/+1*S�����r���TO�\�dM�P��"<ŭ�K���0�y��m`���b+$8od�=�Z1��[�"�vw���ĶmZs����=�i8�Ev\%R�66����Ⱥ���f����]��|���:��w�R�G#��0ي�$?|T���Z%?vw`&F0]E��:���	��!d4��;;�����R��ٗ�7�^�<�6�aa��"r�L�1����,�q�_�i0�WW7��Ci"A��l�:+u�4�j@^E�y���#�z^Y��ZHz��ڵ"���57]z\}�}N���l�@��
r
B�o�6Ymb���)\�^�+����d*x�-C�辄	����=_7�%��94��@Dj��;�;�`W{�
}xE�(��V��Sz�n��N;_F=��2E�o�c͎�s���x7��0,�YY�����V�b$���b�SI<O���]>V���[n	,��b��_�l�2g�7�q��1T�ob� pA7�a�������.��$�&���J��e�T�B$���m!D�WZڒ�5M�a�,�N�CH�7z驚)�Gy��&`}p|���N��7���h<�{S� m_��]{� �*�A_��Sv�܇���D������η�8{�Ն��n��vҶ?F�UX7�O�\%�QҘ2R:�mD�]�u���|!�SF7.��!���[g�Et	
��F=��g�~��Zn⽕4>���^��_��합�HZ�+i$L��0�֭��N����`c�����Vև�Ɯ�hDׄ���>�e������S-��t�j�w��B��dΗ�@P62�=C�<v� ��_����Jg=:B �K5�YNmsn���j��뢐��qN�T��M�I���xT���r��|�s����C�����>���^�6������M@�X�c�n&ն��3��L��Q1���y{���z����QT��OIlH�~��O�=��_>.t*Q��+Ǿi�.�o�]��*]\,�@��	�5Є�u�\�L �~r~L67KN���T�F �0��YW#�
a5j5�	R���f:;�����BV�<L��w���:XD�S��K��ơm����נ�m��Dc�SW�yW9��D
����C�y�!Xӳ��}����Y�㆜HJ�n�;�
V��v�x���K�+��~}??M]����[����J7��Py/.���t`=���v�(�{K�}���j�"�`�olY1���A�4ل�Bd�V f�y��fb��F��]��)�����t�OǞs�"��P�dgFP���)�ەYF��5�Z�ެ��G*��D���V�)��v{���Or�Ȼ���i�5�E�%����k�B�Lt��.�ǡqc:�h�P�%
�`4lȣ�Xvq[��h��O��z�h�%ѱcM���ѝ��@�Ӯzͤ�|�R�4����uo�H�Q�?.�����i1*<���j˘��^����g�X,�a��&�+���T���ܙ#DpPN�@�!FOc��y���69�HOuv�ɮ&���x#Y�WdxæH��l��-cmR��'�[1�T�T܂-�j�]r�_�U��I���*/0gUgu�4n��hI&_iR�P�+v�����5���';��an�"��I��K54�@�J}��e}廞�R|�k7t��a�P��i�DrQN>&x)�� �2=��--ހPM<��_�y����_��b, �J��}8�G�9����K����Xn��%�+]1��4� �|ޞ�?]#&�^c���*� T�8�O�:\�T� ���"��c;	��$���/&��/���I�ݭ�0���6��_�]+���qZ� ����!R��2�㧧�X��̥�x|�e��C��[Ŷ_d��fI�u�����+�]��YR���<ơyr0�p�ד����G�l���b�sv�����������z����O�qK]����2&mV�c�C*�H'
�YL�n�}�����5�E�Q�Ǣ����KxK��$������Ÿ�F�}g_L��@�:}���XQ��5���'��9FY����h�{�z�}/2��b�>O	��kb�����/�Ͽ�tｃ|�A�.(8G���JY^rSb�Q6#B�J)�sx�1�<9�/Hr�W�Z�6f#-e+�_\��z��{�x[�
�(Ƴ�6?�w�P��ч�?�3���_��i3G��Vi�����l[Y���)��f��CH�[|����F3#[���b۲��f�ZT9i�Έ�3M !; �2T�F�<�����y�PAJ�����{n`�N��˙;��&���G-G�i�l	)��7q`���m��H-c,��;9��<�f�_�v_p��|4z�ET��.sY^@����M�uP{>�1r����s�~m�CG�����]�w���^���V鎶XP唳s�d��Iz=c2C����y�Ms}��j���x;@�#QM��+=���f<Q��F�	������g<�sIM��Z�!<.���d��Q����l�yL�`�o���KXcљ(����f"�D�c1\[l�R�Ab�����e[i�~tP��ԅ3���l�¡Vd�aY�kt�oe���I��&M�@, %�-3���-3`0��%F�
��d�����A��'�kX��O�,9O��>�3�`#���L��[-�|hԵ����Bx����~w[ E�ռ�h��0�\d�%ȝ��3Fk��}D�#����r�O2�����o��=u	l9�e�xz�����I5'9��8v+x �ζ�)a@�DL���c�Q��;_[�����8u�@����9.B�X"���l�W��8��z��,�<@���[�,=J2t�:��Nw�@���:g�v�Ñ��͟������A����7�âȐ%���95�p^��(a�S�`��w%���<�=c�u[N\��M������54~"A_�Ԙ���$T�������I!~�<&����� a��ڢp���~��aQGR�
��}*P�Ɋ�e�i�̺J���d�ܹ� ��N��[s-00;��%T�vS1�a:��|�yTf4G��Cy�G[cA����ȁE�+v먐v�:HI.8��t�:�����+��0:R�߽�`l��9Yqp<��Im�h&�C5
����6�YD���;�k�%'�F�vJǞT� �����L�
�=�f�a$�F¤gE8�a'��-�Pb2�3�M ����qsQ:[�H���hB�<�jx���s��e ����!~Y��U�a/~���}5p�������:���Z�AК�~z�H�k�����Ϡ`��M[<O4��V�%�'��1[�l'�|�(Jl?^k���c���H���t�2��;ϐ�g�g�Ѓ��E8�m���������uFÎ��0W�u���g�����G���\*+��q2�5��W���F������3��b�/��Y7�c�B�л�F/(�����ȳ����BnJ��ʶ���Ƙt�"k�h��N23�L��E�edo�ep�(,Tu���5��heSK��NQu	<��z���tq�k����M�� :T9�%0d��J��;$�d���Q��M0����[PEGͻv9���Bl�l<k���f{��?8q��jH+s���$~q� i�~*��IwH(HH�!�X���"�X���q�}MnF�Q��,#%U��CD[K�J�TGIchq��xZi�ǻ�i�$:�����u�gP�|�xdp�J�����_T&�rd�*�!��2?v�]�� 	}ebB"K OR���W�xv�SF��X�k`8�E�L�0�2Sފa'�/D�ۄ�(�J_�Y:��UG�)� T嶡1�3җ�n���_�>���R�a�5�}��V����WH��hp����;Th���������sz���Lǔ�|��q�A9;d�G�zi�fhIV� L��-V]�J@+4�B�ֈR�(b����0Y�LJ�����'�j��,A_���Dr�/�,HZ�@���R�;���b�eeL*s�	�)�͖��B>�_�1�9DI�6��c��7�͡��C���G�R(�:����`��P/G듺h�va�sΘ��CPjN�S��j�'�b�1F��dO����Y�e&��vٳ�4��H��ՕBJwb�ؕ��L�a��뢏�pJi��O�H	 �/���H�)���Ɖ7q�W��+T��Tᥖ�Av(��0 ���d�麰�?}�ҏ6/�2���ZM�#��;gWN1*?.���w�N�ï��ϵ�����I[-�9��əX���`�AK�qs,�>zK��"�˞�aJ�(DmA���y-W�R��*\W"�(��\�u*WZ�C�����n�V `���w����<��}��9���u&G�� <RoT�$U�FL�e�dVr௧L�!A��6�L46�3�* v�!r&I�>�K9��n�<vq�sV��){�u'S�0]x�x��B!����M��x����M���4�1?��z��7朖"�ZbȵM1$����ӧ��	a f;P��tЀ�O��aB|?��!V�m���e��gB@�c����a＇ �N�I��Yԁ6��ʐe�@~��,���fAh�^��b��28��Suߑ_�!�T��SY�Kz��u%K^��_�s��7�WB�m�t��$zde�I��@���<1�J�v�����ԣ��,�}���Go���������죾�s�� �m7����'e����k5��u�T�O�����rLa��a,�h*�Ps�l&������2��F��NUx�ʡ�4h=�8�O��Y�*^#RK6k�G#����2\���eF���c����+0(2﹍�}#�q�=�r(F���K��D!��B�
	�R;U����� iV�����gci���\q�£����C�Mc�Xb��H��\T��/� �"U���◓�2n��%�n/K}�8�Sx����C�+�#t���W��6S���;��[sF��ѓ�;�]��,�)�ճ���������ό��࣠	����2ů^�Gy"��	G���i�Mק}t�DE�3�����e�.8�N`�{������!���=�)p;$��eW��vtvʀ�<T�e%�����=<�ҐbJ��dG`����ޱ���B������|��s�+�R(#q�C�=���^u`L��d�H(ᾡ��BvS��!v��.r���-��
���c\���.TF���(�MFyY��D�����0wF*�5K�k�u���P�� �>o+|~��f�W9�Q�����ey&ÿ�P��Ş.#�U�Bm�[��z�Sj�T`ORMk��脶�m�6��NY����A�j�S�X�XJݻ�Vw@����њ��*[Z��I���瓉��t�=z�P��P�q�ʾ��������j$��>\8>��
���I�R�0b6i�"��<~�i�0/��:F6�=7|�yB@��	�P�Cs�Nmm�Vߧ��_^�
�p�w]��x"H�9H{辱�����C^��}?jљ;�;���� ��1Ful#��Y�1}�����~�O���ډ�{�*	�5N$I�
]ԇ0����?!"���n7��ɺנ�Y�	��D�7���5�'��@+Tp�_��'���ϒ�"��F�^?��j�L�w�����r@-�e���[_
�Z��3'�������!��U
��Z�Z<=��sS�T�D��Y�C���e���ȷt_����ۦ6����8�������:j�ϯs��7J�m��1�}�>4��.�VaE��9�z��w���bFVIyG3�i��91{Dg{g�6{}-� ���j��L(�j�����^�Y��|w{]M:4&T)r���b�_d���U����P�s�K�pʆ#��B�?G"�q��?v+g�${%����"��A�+E�
R'�^��{��gw�m�^>i�v��Y�(&�����uD��aX��f����qS��QG%~%7�>`��6��by�$�j��i�c�l:��v���u��>g;��z�Nk.��/��"f�!\@�C�=�r p�VR-�p���YBK�`h�_�Zq�I�����O�/��'���r���^��~�H~j\���l��5�x� �g7;=�"o�\�QpsaH�x:���P��C�m܁i�9kܶ� ��b!�GX��!� Τc&�y0�Wͬ�R��y���C�Y/�u�J�4�x���}A�tp��m7��)�����$;N��V*Զ.g��Zo�>�s�,�1��7�<�%�����c.a#Ѹ�UA�_'�S���fS�3�W_ȫ�����<,�1̂˪X�����B@��^������2+��9Mv9�<�\
e1̍gV�w7�4�K��F���-y��T���L�!�H�ڵ�c��w}EDX�@���p*��7@�8��zw�����#���&E�fI�,���ώ:	��!t���Zf�#Je�x�E�d�e��^`�Z�m��:g��%��0�*"D� b��9v_7��\�y�W�������������*R@I7� � YV��𞣏pZX����"�w6�w6�6wA�<����whM���#6�T�SZE��wk'��]c{�!���m8�MA�G�y+00���L%;��x,����	w�7��M�[�s����]p�%�w�SS7���ȅ�ޝ�I��=Wm��Fa[�ЙYw���g�q�ҕ� ������������C����g�cb�L��O�X|bX�@���Eު�V�����������>T�9��C
ץ�QK]JI��Ra +x@U�m���|F���F�u��q��s�Tbv���$�ͻ�#\͞~慽�W(��.�t��~{�}Gۛ�+�_�-Z��G�8����`]���r�Ae�m���#M ���D�>�7P�ca�U��h0��	6?� .������&l-۬E�I�(ѤM��/692Rl}[p��m6kp��j����ݞ#;V�}��sX�mHWpH�2�T�K���\J�^j�tj��7�5�Zs#3���'2"��
S��λx&�,�戞8*���7�?mj�����Z^ ���A�)K������<�DIve�K�)��'������N��`@�H�A������'�1��&��oi��8�kB�摪d=@��<@S��X�u�:����m�\q�
އ��+~/��%�C�!t�o� �^�e�7�d�s��{�ja�t���5EhY�z@�sI�ӊ�X~OT���Dh,��5/x��sX|��]���<\X��0���Ǡ�f�P����FJ "z21��C�+(�EM|F����o�f���Q[�w}\H�z3��2�&����]�Nd8�'��F�4r���md&�$q�rc�V�w�:֠C�o|	�	��d��ʹ>�[���Fm�C��V �bЌ������WU��@X��x��37,����>to��F2�H5�l��jW]�|�aa�~.
���a��i܇!W���4Mw���c?���t�֓5��x[w��L���&�R�P�h�1����Hu�r������P�����Vj�g�$*D���峞0�����L���J��D��⚏
4� �c
���吀�Ix_;o4��"=���&מٙc��a��CŨB��WJ�1Ȇg�O����7���R%G��E %Q���z����l����[Vn*P,��@n�8��Α�%4��@��a�����sRh�'�Y5�NCe�]��V�{WPN	׈Bk����ccgXv.O��2>Fm�N�e��4�4᭬3����f���_ϫf���;5κ2�Cw"����m.y�yX�����B;~��ĢY��CK��E{-��c@�0��c"��͂�?��{c����>�T�+S������D0�eU:!��ۆ�uS>a�������9��q3a��,������&ބh���b�<��`���m/���=��-��_�ҝُ�Ȕ��t������QZc��R���:�Zn����g5��1
��C=�t�)pQ�X��'վ���)7L�2�a�Z��#���KN����|BN�wye�2��ԭxe����}��S��k(�u��?;e�a�䤣�������8�tpIi��iHھr�L2<�]+���XO�A������3� .�fi��Z�s�m��G�32Y���OrD�Dg��$�T��"�O�ϭ�,/��B����U,���x���(׹��K���F��N�7��]UA!��  �R(�F���2��6���s�lGkC�i�>��s*��K2�9'I;mS�m��J{��K�=;D��Ol�9�١�`v��N���,F�.����Z~�1�m�݋$��<P�j��
��Q����c��'m��� Wԕ�IŠ�_�����.��e���LPA”���{��K6�)�t��j����N	��_����`F�
� ����}�3���b�:�X�CC��8Q�赯��7<u����δJ.��	�u�k� �!�������T6sR�$�}n(�hKen�RT�?&��� T�3
Y%`/œ�3�$J���'z� ������X���wy}��&�GUNA�@h:M=�S�����kC���#]iW�dc�;b�|�G�
�MB�����^�MV��+a���6F,{�N��(V<����Z늙٤$.1&�c�ꁳ���e�p
�-�C,��D�XX���:�v���b�g7I ��z�uK�u�8O�^��S��/F�N��g,���[�2�0r0h��Rϫ�,�b�ͯ�������3�d�{�D�u��a����K-4�PX�
/j�齁~LA�u��3�'�d�uǝ4�Q��	����M�M����~v�����l%��[��Ζ5J�����W��~I�\*���>^�)�);�q�������襫3_
Q�o��9>I0�K���	[�T��=�V�`�ڴ�w�&f���z��' ..2&�
�[��I��f`eč��V:O���/�\�n<�|pp	BK��q"���O�/C����n�S��n�F,<�0�7���lJ䱊��#)*=�N��TA�@�)bL��Tm���� (�,��USu��=\�s��-1��pYv��ooKi���Ķ!�3Y˷�k\j�׽�)�Z������uښq�BՍn�k�9!L�Z-{e�����,��~9Pnqg�{�M䤊��7�V��c�d�`P�G�)��o�_P��8+��Yu~�e���5�dL_G5�����r�}_���	竇@�k8�L�@P�8fpO/,�*��	sn8��:o��F���SN����y:/��w�.�v�����u��l���%�N��޾֌�ό ��p�#`U6��UShګ�S&ޢ�m�����D��i"Ϛ8�0e͹>y�(`����Q�;�_��,���,��1���t����Rװ���u���SZ):�:,�q5�ǡT���zlo:�KZ��΄���t�Jo3:Dq��@?e�N���5Z�X�Itʲ�&�ǭ�E&���C�f��9��#&tcQ~.�Rx��I"��6���3�:�h�T��ۗ4�}�a�jH'\��ƈ&�_�5��Uu��ɣԈ�{5mV\8�4�=��!VX2��|�4U`����Co���k�7��%z�zJ�xjì`���A�����,-4[�OS�I��	mX�V�l��s���p��:�  �T�?�؃���U���n����k��x��P�5�F:��^��+l������3&y7����c&W��q�����j�&���ǹ�-7�8:,\���G�g;^n��i|��5�J�����+49��a�3�qS�$[�)��lN����_d���m�&�V�[���!�e�"�|,Z	'��`��p)	��~�8e��L~z֘�D_�Yj�k�}�2qEr�GU]��
�$��̶������9�Ed�DQ�P֙L��������W��`Bz���U��r�@B��˹q���v�Q�=9�� D��/Sm�x�P�����n�(�#-� @��|>b9W��`eG���2\��zB-������ա+M�G��y���4Lt�R髤��F�}͖aAC��>9˟HW'��_�?\�/��i�k!KV�c�$�9�bXP8Ro�" $�m���hRL>n���&����1ot97��zѥ��w�Л��iO�VX�4��Ez��M�>�?܉�HoT�^a�|�jL���[r5��6o��XU��	����&�욝I���ˊ@U�:qgo�����رV�>A���)R/`q<�K��Ϫ�j�O�"�d�Lc���[�5>����5�4�m�n�&Ja ��B��3��o�`u@_��{�l�E�"i�5�}��_�$�,�:�3�������NQ����,�|�@��5�H���\Tf�=���j�+�}>"F���V2��\x�#��yzt�g��hfA�8	��M�؝[�1�X�}��������F2ڷ1��d����F+��F� }h�ҁ��ou�Ħ'7
N�]J���������x���j0]9��vG
�����زjn����S#�F"��W_a.��61�Ы1c/��.�~ʓ�!���֪��1�GT�U�ko�l!_�h��C$_%�� U��G��UQ֭�Q���bgo*o��� ��x#bx;ܷB�I/J����#^��� a�L{0�x�!�y�o4�ZY.�#�\�w�\�P�mWa���*&b�U;.Q}r�o�K�
9\�o���l{�QZv�w�8q�T�v	��cous4CK�@{� ���@fV�$�6;�59ײ��ЪT�?�v�غ�TY�T#�V̊??��?�����0�O��0�ʕc�� ��^��Ѩ��4�0�6�/����N$�����A�kK����i���ZO�P� ��X�*(�	0ln ���t�VK����&��O�Y�����ĕ�G�S��򨒽���=�g6Zy��MG�s�~�.o�?�4�8����<@�\b�Ǿg�Sx6R�]� �����~�ʃd��E��DR�^͐�!G��{��>�1F�������p���� ���ܽ�`��j~����{w
��C4Q���q��S��u��]|
��ڏB�u��Vw�d�o��?����6��O~�(!�E���Z LX�W�3 ��wq.���rtC5�V��������������Eל��h����Խq¦#@d�~.o�~�9_ɗ�5	fn�L��$�����Ӊ� bΆҝ ��� ���gU��C2����*V�2�|��o��Ъul��[eɺ{Q���MA��L<2.y�<0�W�2�~+���L*/��K2Q�C�j�I�M�h\'�t,�H	�?�������ϻ��S��w�w�<�=���|�L�sp=	�������AU���,sKV��=���h��y-&�dZI�CFd|����'d�%���� �Ҳ���fv���sŨM���vV)U��P�����5���4��d�P}thqmLY���Ń]�H�6�O��V���t�?|�)�K�<q��*>-�~�0��P�o�z�]Q�w&�z�"������b����+?�eBL覠>`����I�4�
�i���C��Z���Wq.L�2���uz|��u�s?�N�?�X����O�2�� /��	_�A�V
_��3EȊ}d7r�L��;���l⭩AU�I�,2����$�q���Gz�ॄ�F��� v鄆���\ς��P�e멂!&��s�p`f��uMj�x���t���&u>����{��J{��Y�A�y�~�ChC��n�÷K�˲��L�r��cg5�Hs׳�G=�m�7�n�[ Ü�S�SEjWf��|� !=���x3\TI�N��>��n>�z�ےKO���A^"M?���&f+&m�@�ƪ@�L4�0������z�Q`��� ��,W<j֨sF��*����Mք�ǜP��n�<�=A�lYQ��
0��4��4��ծ��=���U��d�	��Ӈn7	����(D�O�W� �q����ܩ��#��zh<�R�3����A>k�D��$�u���i�رZ	�Q�%k��(�CWX�p�CB����wq��f�M�z�P{v �!`8��P t�~�B��b�u�]�]��f�`���Z���D�4V-�3��s�ʁt��l��~� g����R��9���x/���)��D��H�7�Ȫ4ɣЂ���	�I�J���#Л��T�X��t�Vb�Z+�>M)���Ъvh�T%S���>�K��iJ �<�"%��?<{t��"d&LI�޼\�緅7DDF�	���y$`��Z�I�s`�D�P��j�w�%h�B�Kӻ^��<^1*��%�cOLS)׋p������_�F�-��cͨ@&'��	ҚN\���	��b��h&�v��$�p� ��؈{Oq!~$�,�`�*��Ȟ�&`nE��}��|e���#P�Xs�O����Φ<?�c� ��Z��t��(�n]�N�@HWh�o%���`���2�����7��1��G�ey���캠���l�w�#�#oLq�$����9��;�̈́M�՚]t���Wω�K�_�Jݪ�j��"d>W�d���֭ab������a
B'݇w����n��G^�:�\��d�(��D%je:���ߑn�!�>B_s%;./�sJ�-#��&mN.
FW(IW� &,�b�5Eъ��[j�xԊF�x������A�g���N��/�K���W��?�o��d;׺��Y�˥w���R2k�O�Ut�|+����a����f�؞��J��1�#����6��{]���v�>��"�q3&J(˞����	�-��w�C�Q~�|)�weA�2�WxӐ�L����l.�ȁS�
����r	j#N29)��k��Y��k���P�v�~OZ�GI7@^�:�w�S��n�6�x�{� TZIu�dH-Y�+y�c�K�r���|�b�n��.��F*���o��޼�3��J�C	�PM�;�\�<h�F}���R�u|�A�E&��C�e��U*�*֡SW{�ti���&�PԚ�h�
I_�o�\��"Ϋ�������,��/�k���+4�UQ�ã1)�|,@3��`�l��%��*��Ơ0j�G�����"��\�(�����j\�]����f�z�-�(�+v���B�����b���l�a�,�ϟ1���93D�z1��H�*
���n��W��.��Lx́_a��|��a���]ӿf�|�3�=$ꀲ��A	k�JC�8�*{-{DP��\م�
?�^<��Ⱦ ��W_D&z���Î�?EB��N���> �4Ԅƫ~$sO�]� �A
خ>p��АI���l���dE�1!�U�[�j\zԢ��c�J��?�S��wwyv�^w�Ͳ�^�����Ѫ�p?E:��D��ZԲ�6酖��M����'R�e�[\n���ζ!ukK�B���ާ^���c����~�.s�Ҏ�`��DhI���!;/�ߦU۩����Ũa�e&q��+;��w��يTV�|TW|�_��66O�ʰ�e'��b�Y�O�=�E\���#I\�(m<R2�qH���s1�Ҕ����+����E�=�'.�sr�;�zp���û@�©h�� |q�+��L���->Y=;��e�����^V��`C����C��e�H�&<QH�Z�ۜ���"!iL=�����L�s@W������c�ב�9Ւ����C��$�v0�۾.hJ5j��&�ڴ�c�\Qe|`+o2� }G�}{�,��S?c̯������͕򶨚�Y�`�E>�{�ۧr3��7�峴�|~��N�[���׬J���)mO�' ���I`��e _�Jg�a�0j���%(!D�n����x�d��q|��Q\��8v�rݝۇXƵ�P�U3���	/��*�i7fm �l��ʿAj�����b�2�{w%��B���dUwdM`�8�i:�+�;���؂݃�G�
�iw^��e-p�@��V�����sW���<�ɚ{LIO9Z�=?�W@!�FᩊZ�������n����V����/�	v�����R?V��Џl��Il�!HD�sXo�����';�h�˓�Ae0}r��c!}�W�[�����
����*��(��@�g6����C�`@��y�� ���.YÎ�T��"s|4k�Ƽo(���	Y�~��k�&p�f"��l��٥&�2Q�Ĝ>���zE��k�W�W�2������/$m��l��D#yw�U�A�]��T\�\�اÑ�h��db�U��p������:�+V��g?Mi~V̮Y4���o��ծڟ���%Y�����{�h�h��N����#"Mk�ق i�H����N,\�r�������V����x����ڝ���vN���
R%R���L ^���#�:͸�;t�H�g�\w":+T��î�T��m�%�o�	���w��[4Xu7�r���k^�w�����9��A��e���}�\x)��] x��6^�)�<���|�����| ����?^��?Ѥ*G�xQ|�*�_�p��6���U�>�JQ��(�%�����ғ�l��(��;�����.�m�ג2��>1��(����9.���5R<���%t������ij,M���LJZ³N��2f�S�&�(MД�y�yI>�����*�������ˤ-eL�_��B^~��p��Hq����6FȰr/g=�K�N�͞x�L���F|�GďDW|(3��߸C��mM�ϓc�+k���N���b�7�/�9�i#�
�XF#��P��t�A~!�S̯�G_a�&�,�>g�'D�C�U�6��%`?F�_>��#U�Uc'�L��l��/��K��y�9��	8����颤�B���G��4k�+'�#�)�[�8�ۘ��{\0/�j~��-�b;HN'�%Uq�ɭ�O���tJ�/^
����e��82�6�]FMp8Q�A�5DY��:�4\t$����$N�SBHxN� L����W)�������:w0�[�m9�xϙ��~�9�D��aϔ+4�2�x8<�n�|����R)Yf7f/�&�OA�N�=k>K�^A+�n@���������mX��#�FoYQS?`����Ҭ����|�����n��P���M�]���_�|C�4G����˖��T9��e�-����x8}�� J�r��#�;?�Wl�`q�q"�h��O�<oR鎘'�f�����Q�'N�'�BБdJ����v�=$��T�&k1wmk�shU��t�m�XK=���eΥ+��1{0E����"�â�H;�����ѓs�$%f糸|r3�B�S"xa��T�*,~��H�%C@Uo����4�F����1+-rЂ�9���6A�y�]`��Iz�!�]ǖ+����ky�;��ϻ���)��B�ѮJ��9N^���.IX�=� ��G��I� G�>��J�~�Wg�С���>ˣ�Az��7��]:U-���x�E䋞���$ޡc4�������q�����2OSԹ8�d��p.Q��<��|���*��ߚ��}yv�ϑ)MC���D��i��蠦r�XW,�S:�0_����PB*���/�_>�$�����G�ͼz�K�ŜY�����s���e��Y��v`�%��ٴ�� �J��D@��5�e�W?1iʕ$̨�|�!M�%o���@te��óSu_:�:�7W�m=�j��@6���U
��k�|�M�L(�x�E0�uP�����}���J�{�ُ]�k��~���ݴ>���4)���[�̕.[�'�?�Q��$WH��H"�X�g �t6h4T�%��ga���:t_?��Z��Պ��8��5"�)�-��M���q�V�E����Ϊ�;�rH�{��m�K:�H������	����|�%a<�#�#���]g}S�Y�o�p�ܠp�>?�hﶋ?kl|�=��z��OA�!\��	����r��@��� v	���6��P�	��f����L���x�*��OJ3[e�"I8�ڀF�)���r�R��P���S�`�)K]��lAPA��aE���
|a C1S��!F�u��iV Y�_U� zOt\8�vc��D�yS^,���+�_J'����e٘�)<��4��l��4���K��ʘ_�]Cn�#W�^~��M657҅�E����)<��֖V�Z7QE��%_C0�Y2��9���F,)�3�d���y2HPZ�YJ2 i ��"�}�q�`�F��گ&N�F	`0^��`��v�G�L�\����	(9u�Ղk�Ҕ�o�r'"D�p��{/ì�@j"͸E4�<lpza9p�b��;h����<��]�N���*"�7(��� Nji63U�+�[�ŵLE0� J��.�-@Z���@�n�*�����y�N��y
�_�Ӳ�m�x>1Urٰ*1u�Σ!��v ������N�?G�`��	��a�7W�ݍ�W@㸍���IҔ=�ғ�|��Pڎ�+�mh�0���{?J�Y�L�I �S��:���a��͒>�#�s�%<�hs��H�jb�$��p*�m牍���N�;>�ƙŤs��-�5Lh�[�Ŀط��coP��}�럋J�5���4<�P;��S'Ln�rW���P�.�ʔa�ד�M}�َ�d=ܢ��<���7Ξ�N�Y���؅����@T����7MW'��E����1����6�k�u]�> j�my����2��垾tw ��6�����<S%M�qN7��+:���AP<�{]HX^�|8�wQȌ�������MІ�B�.H�}��Jd�@B�����/��)�Lk�u���o%�J�}���Q���m&R�z)�TL��t<N�}��D~�w�$��n��7D�(�r��5������)B����:Փ�zo]��>���wB|�ڠ��~���[��I=<N�� 6��z�~�P�����0`;$��f&�C
G[qd�K>K��"'g�a��v"%��@?��A�IE&$��Q�1[L�f�������U\R����i�W����8T'�r�?w�t�L[&�5���V���v���t�񳩶�;~�Ǡ���@�G���
�K�zi#�y��<�?�J-�=�����:�"�y��h�R��|��j�s��=Q�l�'�̅�ս�H'��铍����ʈAI(f��m�����/J�Zo��P�7y�s~a{Ц�7ʌchK�R`�I�Q=�0���='y8R�E#C8�8pQ�q ���w�Է0u.���F;��#�j�j��q�7�uX<�>�w�����~"(���^�|��2�g;��ɯ���:-o=:TV �����U�w�؎z�F<~K�(�l8�n,�Mmhԃ�x�o�����Sh���!��z$�]�b�!�	���cBl��i:N�/�)�����e���񎌫c��x��P{6�=7� �8u�s ����	�{�ޜ-�����K��Нs��C�U�XΡ�{�e������0[[�������S������C�w�PL�� �:N�ڟc�eG�w�{��������Ov���{���+���yy���6�2��Eh�f���@i�xp�G��;�A,	�����,5�;W���Xz�ɘiJc8i�0:ܱ��X��~��bI6�o�;�'+,���5�O$j�F�yu�#q\'���B��O?����z9/���;��wpi�T�)��ޥF���ǅ�y��ո�/0h�79�RA�%��O�
�M�N����öN�}�؅$��ٚ�C����N���Р�xaR&�ïP[��E o��J����d.YV����<Gψ99ʹbᇎo�d'Y��A�vXR��x�n�D6C�b�ܶ�y%��խ��v�|u9�T�a��Ck67���xÎO��we��~c�SuTI�/B�8�YƗ�'�[H�=~�f����[���LAX�ՈKh���\�>�q��*��I`���D�ىe����b枎�$�꛲�^@�Kk�/�[Rg�,�q,��At���J�lݳ�N��ZO"I"S�7�S�e
(�z�%�I?9x����Fu7ez
GS�e�Xc/�X���J�OA�^�u��==:�_T }���%V�R��C�+?I���%溧//�ew���^
����$������QI}68�}2l7��G�uZ����2߿+X����D�xT�-�Ď��i�[����gg��|7T;O��e�7�?{uӉv�*k�b��)�?�0g��G(�ۚ.$�a��/qB0|���R����'�5��1�ͤ�28ueiL_1�J�yb��Ȕ." ����H�����WL��0�n��8�n1)���}Ǆ%��&ü͔�K��d;�K��D��bړt� 3ռ��Gi1���6�
�e�p�UhWV��F��`�z���{BK~Gź�|u�7sE�m����L�̑�0��-���r' �數<�>:���Z45.9�Y}0:50�����U�i\�v�?|y�Z�&n�*�8��1+�C�a��~�j�.�e��u����mȏ{t�R?c9��*�St&���P�2`�X�Q��݀� ��#+&�bl�t2�����)u����%��r�v�d�_	�{����D�n9�8�9ơ��Jڳr�!������'��g����߿u`��F�;����"��e'�h�d��N��+�S']��f�ڀ����ŷ�Ќu�_��]yF��=�����w�W��m�C�����Pt5�f�lR�v�77(_�e}K>����Ķ�g@����\���7�<l#"B2�ZD�r�@�J�-d�H����G�qO2�D�.�b�M>�g�z/�s�p�����Fĭ(��H&�si�,��ej[���#r���(�x�vr˥I��	DO~�o�բK_/�~�V�T/d�H&V
3X|��X�n�	��^
j��:�rH�n��ZJ�O�e����8�<���}�t�����+j(~�i����?����ٟ�k���Vϳ�$�O(�9P*c����>�|B���k�vrCPV2��	p$	ީ�B5�[���� ��L�o��O�ڶ�� [fO��L	i9
Jj�S�їl�~MM�Pb$s�Pr�ŝ#ЎA�Ŗ�_��5,�r�BJߒs��8�lW���T����Ch�PɢK�pc"9'��S�e6�♲ᓜ�(�yZ�+Ӏ�օO�s��`5�LW8m�)�I���7q��2=��LRct)Q�պ��OuTj��tP�e]��5���K�Z7M���KF�ߚz��w�đ:�|�#96��[�ͧ~w��F�R��}�X9M'2�lgQ�Q��S�f�ַ�Li���y��2�l�xL��Bv�ɾ�Mם���@HQ2�b��"5�����Ѐ�����7#�G���}�]6�i`琢��2�yI�J����&~A>���_{����_����P�[p_,#y�a%}*1?kWB�Xe�έu��#Lج���s+�l�Bi�l�1;�2r�A.�ؔN��,��E�9Ă+�l�~l�)����\�z��7Ͻ���E��E�����!����3/��r6w��M�3��e�\N�������jh��#{dLx����Z�K��ScK�&�����5��`��U�z�A�dC���-���.RH*�nK�*��/:�L�����1#-F�b�,~O�������ۛ#����|͙)���O} ��O��3M�cOôu T>O�a�y�}=bP�֟&��/͟I��bيĨ�b����C��l�Rk.��	ź<��$K!L���K�<��/���2%R+�9��+��Kډ�w�+H��ghw�Cx��%�n�M�nk/�
텤i�L����:TIFM�)��N�^�3�h�a�P�)t�#܁�(�M%���o55��q3����ϐ���"�0�٩NA�c�s�0^���j�)�|�m�=��<�.곦d�W��ܯH<g��#�ҡ�y/���c�U�V�PCo$#��'�Cw�缹v��ێ]�jʧV��D���f����ؒ�d5��XwT	���(�*.l�G2.�φ�������+3���~++��M�-y�U� ���y�"@�OU��f�Tn�2y�C��J`2�?�{�TF�Ze#ԂN��=W��;m��Esg1������E>�M�[lS�&p�x~�����8M�2Ц)af�l� ޮ8���Y�te�!�	N��ހ�l^�~�BV^H�������b�Ӏ0p�C`��C}x�@�[�<+*��N���Q�I��;����XD�q%O��I;	ٖ�i��R 'F���=���3_*��y��HS򛎕3��!��R,�P�}v��av�^ݶ._Ҋ
���s�"�,��D��� ��;d�����OA�Obq R�)^�خ��Ң��h3 E7�/*�|b�F�_\��Z����i1u|�d�7#@�P��L
��$��v<�D�^�VgҞۓ���,���Fs���ϻ�:�_�_�Q���h�w싷\�&��r�G�r�萲�UM���ߥf�^LI����I��%�8t�s(��׶6���T��O��ğ����+�`#b�$C�Ǹ��	���3%�ų�n�4/�bnB@۵��G	��y"6\�tvh���bQ(�,hL*�<>*�*�5g�g���R�O����J��I6���@ז?���"�5�<uAms}��X�d�O>���t�1����`�dH�7�a�;�:����)"�I��3��I�-��L��``��ui�r*|+��|<������Ѷ`��"�T"���! ���;*Rӿ#��,��V'��:j��a�~�JB\�U�C� d�ݔ���b,��Q�c��Gfa("Ey����:���K������m�۸�S�Wl^3ƢH�:EpRR����L\�Չ�3Or��P�]Wɜ���}y��)6K$��Z�i�`g��)�5>�?�a<P�y�s��O�%�;Ez�>!DM=u-*��W�w�b(÷��4�e�`�*1�6H���c�p�,e����B1��bn�s�ѯ;ȯ��O��k#�||�E��j�~>�O@�ϓ�U��i��_��������u�8�#Z�R/�Eo6q��ŧe'�]��@�f
��xC�u@�?�}l�{�V�O�Ԫ�üۃ��%���ܦ=������g;�#y�F(�L	����R�[�qt{{�{AO�:���.g��RJ��\5D���2ch?�l�=�<�+JĀ����;4�1%d�$�g |S�Р��*C�$<V�h��c���O䇖t�'w�e:.���bͲE���VAH}i	L|��|�7�a�5q�� R�� ŷ��'p���%
/d�St%��q�Й�5����.�.&I
˫��Oe�]C��y��ުl�g���~ytK���ѿ�H%�4���A�a�-��N#�Ϟ�+��(6�)���n�"�0M(��?���O��f	h�����l=.&k�+UlS�C٪�IJ�9�u��<oUoh\+�|��iL#��&/|U{��݆�N��e����* M�8H5����w�2�L~�Pd#kK%t���&[k���/w����A|Ĵ����p{�m��h� ���F�����iº�W�~�mI�O�%�g��\z��ඍaA��L"��hu�Y6��p�  ���Y)�l�c��jA��E`�\�7O��w��8�˅OT���-�Г�B_����G3�:�~�F�v �9�*��b���E\h�U/@�4V��o��� ��%';�����ǩw��4EW�-?�9>Ûդ}G�:�ݿl�<�A����Cb���������0�Oн�$�Wo~�8pc��D��HR�B"`?�t�ܙ�ǰs�^Z��	�H��X�
�F�q���(ޑ%���a-��� �J��3�c���&L�� ���Уr&�3�2�]�q]/=ߌ�D�I��Y��4����)�N��_r|[���D͞�"Q�%ki�kZ0�<�(q�ݥ%�c�'���0�rv�:#���Z����Q#��9�����XD8[牲_dk�e�:�ޡ�"�e�g;o��'�d�^�S����o��_�Z�w՘r��\K�v�2��ǽ+�T�Y-N�:��	]��1��`*/�v
Mf��^��~TJ8�Np���A�X8��:o+S&�%��u,��{�z�d#��	��cԱоP��Ͽ��ozo�t�\W��)�@~ڥ���tHw#�J�U��
�/���u�Ub��,r�sĒ�i�4��s]Z�[��ͻ�U;��A�B��b/��*�)����.ު���0�q��(evM�-ؘW�O>�I�V�N`�]pص�X%?�V?�߻��M|x$��5����1�����x��������kPh+��`�(�[�*�
��.*P�� Ǫ�q���^I�� �eT��䰘n�5g&.K�YA%nH���?���VI��@A��z�����9ڹP(�J�H����h%@�xdk�9Rr�_�t�"R(���O�Ń�A�41EI�^�|Y�������J��-��5pP=Vm�c[ނȯ��D_���%��G�Il� 	l;̎<�:�O�ĵ%�d�+[���O�i�MB���{��c� u��5�qJ�����Ҭ�ojx�{�V�)*��N�:����i.�F�����$����L�!P�o�8�xW(g{��dd�;EP ��+Wyy?�����g��/��#R�`r��?�����Y��bs���)�L>Z�gSn?��q��5f�5����$l}U�G\ul�YT0'Vr$�q�c�BË�Y6����ʊ6쥫&p�)Rk0Vx���pX{������E��G�1!�2)�9wVe�:�kv��O�g��7Q�Q���y�X��lO�)�ُ�g�Dݝ��*$��G�Zf�7��e�������� ٰφ��rȜ�1���5}vV�i�P.^Z�0���FG��R7�Ւ�M���0�c�}��Z�o��_�����r�%E�ow~���|/��ǝ6����b(�k��co%Nf��K��C��{��۟�W�=[���Ňl��GWܴU8c�0hMK�>	1l��%��]�M�f� ���Y������oHL�Y'K8ĉΝ�<�m����z�\َu8�R:v�����:&������S1LV�j�CqS�����`Z�~���7G�|էL �c\�����6�Ck��o�YQ�JI, �i�N�r(�/��W�M������YQd	���)�?.z�^�	?��u;|Ϯ�u�~�գY-���b*��M�G�sQ��#�s��E�"�Ja�8�ƅ0/�ۖ�|$��=l��s��Ҙ�V�SWi@mO�oN�<�<NĹ�^�8����C�4�ü�j��a|EoO.e�@���v�mr���p�˴��@��1��h�Tu���mƍ��$b��zj����@��)��-��A+��X��K렜[i��o)*�l�|m�R����<��|��/"�.����$<Yr���
��Y��B�C��_lO�I�5��}�W��`����xQ/b��-�L_�:������?�.ʆ����o���g�i�4�Xs��3��B����}҂{��$#�h��13 ��1�����m�a\�<��5g�1�Xb:2����:kx�i��P�)^]��$h�[��E�x��g+]J��i�����uo3�9�ի
rt�H9$����=��Fc�|J��!�g�_A�	�|��8?�V�ʰ؛�'Q{�T���]5}4D�����u�x�/���X��=<#.�|2}!�9���z�,^ϥ�N�����DG�_����x])Ƿ���]Xd_��sT��ﳇ6�b�F���F]9� �g�h��(�G��`�Z�y�F6]| _�I�f�S^�f��}��g���e�H^���WmʈZ�@#t-W �lʠ���2ʖ-��ɜ��VŇ�
���,a[��K��܆�ٟ�8m=�/r�L�x���W����E��0j����j8�m�`��툦���l�Ê��ÉV sZi�U��%�|�y��a۠�>b��w@Q�ƨ��5d��7�N?`�E�ۡ�ύ��
$y&�'�#O�����Z�	�����D�0Q�"o�fSi��x�JP6��]��>MX��tet�\'�*��H�_��V�`�s��� r�	�ȑV��ؘ�)�F��k���Vw��%���Ӷ�tI��Յ��x�7h����Nimq�y	�{�K/��
p4�L7���	�z^��Ӄ��W��=;���DVA�0J �����:(mx��݋`��O�6�ñ��x��Ky95h�)��me�,��dǬu���� ���9�:�P; ��1�lK��A;:��O�Y��/�V!%姂��?q[�vlY��$��.���)h�>x,�o��w-13�R���)2H�ms�-�;�o�Wh ��O�e�H�s%D���c��;����s��1�y�"�,DH_��Q�P�=�����k�B�n�G��a�����샧*��5~H��^_@ո�l@Ơ_4z���t�'���T��p���}�Z�>}�4���b O���gz7<�v	$��Rػ�L�C�X=׳�0��I���B $��������
�9 �!�j����e��?uf��VzQ%��$�<o�uز�]�S4�������I�����ܯ듶�?F쑶qR$@l���80�\�ӫ�<4ޢCW��H����.�(�cl"�Y'�+��;��,8Tӽ�kN�=Qk�u��Gm�(�N�+�R�c�2�:x�z
����n3�;�/=����r4�)��Q�B�ԍ�o��d�|uj�u�!	�^�2e
��Y�[]I�Ӡ��k���^�͎�_Rn�3��`�i�����/O���kI!炯R��Yp�Q!윌���cA��
���GzL�}�i���W^=^�}�4�BϜ��gT]z��mrӃ�Pb(�
�S����3�����W�t�䞢����RS{G���D�@f����P0M�2&ք�]3�yV�#�/
B� �}�E�_�L~c�P
m���P� zVN���r<�5C ||����L�,��rX����Z��`�ݵ�g�)�X���l�*�������{j͆&��j�H�N�Rf {Ks6ُ2u����Y�)|LP߄/,Y�J���$�����"�J8�4��s@�e��d��̏�bނBa&�J�T$����W�Q�������D��)d7������Z��b�m��y����8�`��Xt�@N���;]5b�匀S��ֿ���m9�'�N�`�y͊$�j��p���l�踰�@�;�[���7���ro�;����^MO�1=��On��"���%ԝ�`pZd�.����{S��ܬ 6l+ ��Ī*b[��r�ҩ�Y��A�{��-��47I�(��[{�u�2�L�{D�M�����/q�i���ep�����e�����Ift�1xS[Y=���k�=�n�Mv�U�h��"a\�P���%I�⤑v�����êqG���������v<پ\�ӻ]���p�9ox3	O����p��J��p�V�Ȳ�$�eU�Y@����8�t�wB}��ń�th���'��3����(��h1��ڑ3��#�*��ݔ��4����EG��.j*�=`�S�[�VRf�V�����ϑ�d��U�ʷ���*d�q���Q2@����+[���#��/�%�*�I�-|�c&����'��J��D ��ێE�y���>8e�)��{�6I�s�7�J�P|�vɫ�/�BM�RՊ�4J����E)�_E��@�A@Y���T�Cҋ��Q^�rk{,x«L�RbL� ��]� ��7����e��������r��3�	�o�{oQKu�Y�s���{��ZI�;�Y�]�%�gbWd5:��ow�����ҽ�J��DOr��(�J�{�0d�ߋb*��~�����f��KS��HI'v��8�2����*>@m��\�Y�ז�X���5Y}խ��7���D'��_ٵ2�n�zU������-/Η!JNK^yW�m,��7��'9)��Cp�������x_�"GL�#�����z|{�Xj����K!�'�Ր޽��n�[�iJ`���9y�D���.��7,-n0y��3��M��}��q�b�{�C�f�t��������u��ە�fq���I8$�v��� VWAgf�hj��][#ի�,m��5���I2Dty:�l�����Ză��4�b�+�"��X�rP��&7�˲J��_�k��WZSq�mJ�}�M�2g�����L��.�Ql�+���E|	����}���0���f>�7���oC��t"U�h�8	yf�d{|R�aY�C��I|��ePw��h�<�K���o�{����L
����Y;��.���y�uE����9K�ܿ���B�����Y��p��k ��f����e�������t��&�a��(^�5�l�����kx9/q�+f�v;kk^GW����c�#��Q0#��%vR{h7&�SQ�p)����6F���	\���U��!z&'��RcԦTa/���}�6��L�?�a�Z�2�m��6;�Q$�1}k@%���&p����/棓�q1�z�qX��"��,N�v�F����ԉ���_ �:�Mi\�j��{�!z���)�8�F[�M � ��I�P+N�.D��3�?��dI��[��	o�,K��ul 9�6�7N��6#UX^��:M��6�eG%���dp��˱$�c�=�B�4^�qW��Z�*B�Ѻ��j.Ya���t��Y���%��b�ϣ&#ԝ�l�ٽw��Ct�w�$��`}�(���X�!xs�=��s%���!�Z�tK��tG)�D�Ԑ����[9F4���J�քE���l���}��h���0>ŏ�m�3�$5�s�o	ىă
m �Do5����\���S^�����8�8���k0"z�r�[wx��t�ő%�o�Ŕ�f&��؜J���>�����V��M�����$���%�uv��=%yt'�@iE�,��n��[�[�W^؛�K��Ą�������G��G�V/����̚��V�0�K#��� ���$Ǳj��td+��J�t�itDqd�Lf�C�o��n_��q�4���O�9,b�6N�I��z��+��a ���g�7%"ר�rN#Ϸs�6M�~��ٝ-VI�����-p���n�=�����[ #k�x5�����>ANć7��/�fD�&��r��(no1�K���>�j$�_�4U�!�?k���}Ԯ�Fr� �d� �ɜ��n�E?��y+�X��.�(��c*��Y0�Є�r�y)9�����݂�qF��ǿ�O7;�}2G\'��J6Lc��s؎*���%��M����
5�"}&���YZHy���PQ0]������/�ʀ���	C�o�A��^"���4<�+=n�~Y�Q��M"���h8���(Y�hN�ε��N��6b��k���^9�����\	V@�Tx���B�r�V~���7�)�>{y3sKc7`6O���ݲ�͖��<��8G��z�����*�r��kY���� vZP>O8��]���"����� �y���LF�����O;Ԅ���,��+	��}���氠7�V���O� 6��UE(�
c���!u�� ~8�đS�WN�-���*Q�9>����/�aIϒX�;ެL����vK\h��z�a0�Yj⫫ H`������t"������T�I���#Y��Cʠ�ͧ�C&	�}W|<*<������� "�̃�(_S�J�\�[��a���D}/��5SB�e�[裱kn�f��E6d���
����J4��	
�2�	l���FdJ ��X;[N�R71_�n��v��$P{i�R��'Î�[^�����0���0�U��Ш�9��-Tnp
2���iJ�iP�j'O��n�-m�$8l���2[��E턆`?~$��t}�X��:��$����,�uh��lb)�
/{�Fق��AE �Ga�:jgݼ���)��&U�'����Ry.ՂO���>Z�'�5-}|	M�
AZ��шY�w��GvÍw�[=��8�&����y�twQ�{�q�
%�H�ƽ�)�A
�ݾ�i��a��ǽ�Lk^aR��,����&Q�%Qq�:ԕ��绎#�c����^H�~����ʰ�Tm�~z���*���v��놌��U�S�p�(
]����$��Y� BY�h�����]�H$b����ګC'��F0���곏���G��~�XY�(���o� �D��n+R`�8�jī�5T�ئK�&�i�/\��<�������S�/��gH|t�L�o{�C�%4He��f���q.�_��&�&sF�rg��{�D`��I9��zo�ɾ�f�z=�*�x��b��n��8��l�|�N�5L��7}��yH"
f|��ZC�\ہz
w�L��0K�X�;s��3��?7Ǔ�v\hi/b&>�y��A���?�*rg���I�V���zq���3�˖��[�&~�/��\M�(�7�e-�;v���q3v�8ܑl�r_�-P	���˪��E�.�|0����!��d�+�i>w�,����Ě�|�?�����L97����g|�A�����	@�DC#$��\B�>��4�2��q���鬿qrI,[�'���C�&Ʉ 1�&�g�����Z,��6�X�Hyc�ZA��+{����_��K��/O���C�ə�d���") Z��\�pz]�uH�5��t�*��~��淼h�	��S6��/Z˘�u:���I�K��`2vx{N��Rh�"�ȕ�/�n3ׅ���`Xw�0���c��a�l�.X�q�bm�̑D9X�m�-��:NH��,bf����ǉ�'9w1��͑PIi�g�&��[!Y(r�>����@zs�/F�0�1�N�.n����v�t�ß\9�6�]���U�&3j�@g�+���6�z������hP)	|w.&��n�[�e����c�ye��?
��ie�1�����o��Զ���¾�xZ,Qc�f�Ǹ����Ԫ���C�xh��0^ss��ĳ�����]=O��+;e]OlA> �?�)İ.`�]��S/�����FS�r�ٰ�<�;%���M	�j�,)��X�e�J��:3����J �Z���M;g���$������3��d�R�/U.�Mb4�z�A��M�g	�0C���r�UȐI#��m�&{5�A�5z��S
'�m�\+t��$��)��1-�M�u�Y�%�:q��p��' sM7�Pݜ�ճUc�<�q�GN�Ҷ���[Z3��[Z��V!'BE���켄TA÷�v����vҙ�����}�?��>c k×�Kp�#_�ufnS���Vy��)pj��]�䋁����v��%{><�向=�Z!aqa��mGM�Qq�
|`.�?�uMt��P�2W�|��i�:>�g�-.u��D�Q�w�9C�K:�x#�9�,mJ�_f3�^oinT��:�X̂h7�H8y�J"	w�kt��"����� ˓�[aq!�[�CǊv
q�(W��`{��q"T<��=����6(Z�<'?��;�#���6�������	}��V�0�I�����W����G`��ð�a�ސbJ:�'l+����"#���+ō�u�#B�u��o?�٦�R�M�Q)�����7+�ʼc̊��^ľ�B)��hvʌ��u���X
��u#��T�"���0�ǎ�GG�nJ�P�y@�O�b�YثѰh����E�|ZZD�}^�{]Z�|������nȤ:a"Ra�bˬ�>��{����'���`[z��8Ws �����W���6f���s�)%��ﲊ�i� ��ƚeNI>/vh Z��X�j���f�h� ����
�Y;E%���s� ��D�M�`�ʂ�O�ܨ+Z�w��3���A���W�H�X�k��1�5�吋O����[���=� �p�b� Y [�s�@{v��0����K"9!*�4sc�q�C!�qua���伻F���}v.���J����ޢ,�ɥ++ם����7$��ƚ{<�6
	=��8�jn�m;�^�o~:#��Y����T��A.P����By�_��>=���G�꾟	��+��w�8�΃:j0k�Sd�3W$թ�U���(f�L(�-m�`Vєx(��i�OpG�ށ��� k��SQ�3�&=I�,�,��3U��H
cǽ+iW\��7C�p�jb]����Zc26��<��pH'�XGw;+ߢ0��#�,2bn�g��5�U-���n(߇P���[3`J�ri�%�V<f�B���d����:b�	iv�p��9�{}�AG�U��]9��Q<33��ь ^�g8���!7���bJPɺ�(�@hyR4���:��r+T��!z���E�[�=���j~�>-�MUEi�Np�x��Ϊ�~iR�]��!T�E$
m��<\�w��b�_����}�*+��W����,̠'�����a\�=�<׌�Jǜ���-��/�ݑ��� ��a9�����[��F8�d�*è����	�6�rf)�c����d�.���-�CMSwLE,)��+��c�D+�h�2#�٠��A����� ��a.����R���k�/{`���/�,��8'ޖc�T��M�j���>�Z���p��a@����L���"~ pCPI��T���w��H�8Z���8�,�j�­(�m}�tÐõ���̳�b�w�ܫ�;>X�I�s��s�����#�����,M�b�&V�]�'`���Hm�7݌�����P""�W�q��qBh�M�5����
��@���zq�d?���Ţ�=�t�g#����gc���G�O��ڛ���^�۠l���,^[i��IxB�o�N�#n�O`!亅��#3�.4��:�gEO��?�3�uH��5�N)�a����<Y������!�����e� /:]IO�Gz�F�9*}>Y���xi�2z�v���j�l�3��Y��0�����J�ط���}
�K^�̜��P>>[U��Jq���@�K\ۍF6���©���9����J5�S\�`oy�q/�M#�� �7lE+o�f'9�E����+�*ɼ����蘐��^�jU�ݪY`ＷpM./�N�+�ĳb��u}�ȷ�S����=�eѮ{�Q�)W0I��#�Fj�/X���>j���Ĳ��mU�Qk��'����b`����r?�����Ll�0,�v	�w}F4��l�s���)��Sڕ��V���ᯐ��n���z5��2~Z�;a9����3\,�&k���9��
E-Jr6�ʽG��8D_�c�.���vXdg��;�o�	�f��]�Y;e�)Lώ8���@��[�2�46'�Od��ls�i@!�v,�1}��qc����.�#�����ń��D��ބ(ĩ��Rh���t��&��%X@���tF�d_�ls���%�;<&64'�;�}Q���,}:b��Ԏ5[|� ���a�ʤ�Y��2��n� ���}TXv ��ϫ��B�%���$���~m��U��������$	RA���:�o9m>��n�/*E�u>"�~�(6O��
�w.��k�8ɏ-�=S\%f�������_V��R�&E�QXC�Jr���o�8R����^N"��][�}�du�8�w]�r��(���]4
,�\�� ���t���B��du�G�GG#(���Z(覎�DC{�ŕ!��ـ��^�ꌗx4@\e9D\�x�l�ΌWc�0�j���2kfl@�\����:�i#��X1-�(�F-؅�N	��<`n����i�W�,
�r�mLr��n�)���N�Dn!� ���]LE�1�8eG%�L��a��#w�2P�!#&�� �//֖����@n߲oY�6}��
����}�'���4���瘚*�$���l���?#���M��J���֥�J��m�_�<����]p��qk�L���
��:L�x���&�{mFA��������u�#	���8���X��+)1�f�)߱x��2G�\�E].���MF$��Z@���H�\�^���ߵZTX���)>:t0܆H�*��xG8����M�.�Hx!�������"92�'�Nd4"�S�v�n���ɫ��I��E��b�5���W�t (�߳�N��_�������_�>9���I,�
`V�k(���}�?Qƥd*c��6�}$/݆Q�����(�T�{W�&��Ֆ�Փ+�w�H���á���n����J8~��5ȐFO����~Սٵ�َ
�0�#�I5nƜ�sf$8w:�N^afQ�9	��w%��:�\�\G���
xW4��@���Ȓà�do�x�e�Lf����@�̜2A��Y��RlH\8Rx3��Ge�,�KwX��`��&�W&�ſ�4S����/�'<��Q����{%;3��L�Q"}Eq��� ��V�^��_ju])�:f^���Ε�{�{���obD��;8�������ww���N=�D;�uZ�u�\�Au]�E#��d��6!E���|�F`W��W޺�q�f��An���t�1{5$�w�\��T���$\M.�5?�!���p�Y1�A[�3zQ�o��̲\�&&!:�u�~�ݧrZ�ߴ�;�<�s��`d3a��VV����.�1!���KD���:�B���J�&�)�?-nA��/����؆I��p�+�YS�' �vI��(,�s���?�#9]��ZU'_[h܃f5@T��\�
.��b9C�w:�pg�;q �қ�,2l�~�����@a��/��^�,�l�Q[O�%��/�/btVR��h��v �uh��.ـ�`ڮ�'�}�� lpW�j+Z�lp�/��~7�;��#�*�3!�f�|�ضC��^���𱴛�o� Z����1�x��!m�x�8�%���F7�Ay�I({�������?�L�5���(pV�%���𛂬�j�(��Һ�E!�'T�(c��I�m䷢q�b���\�<߁8������"u�؈s9��St���'�t���_} !��rj!(�v"r���ޭc$���[K	�ϐ��#�*}t#\��-a|�B/�����j�7����xN��W�@�t�3{��sli�=�>�c��lR`iH!l6�vb�t���ə��a@���^��A�6i:�L��"�SX�F�<�o���o	�ok����_��SK��jͶK�I_��_:��C��ǿ�H��s��&�V{N��ZH����!ӭ�sS�G�bN�^��0H�������gΉ�,���E����$.�,?��kB��dĹ�aU���؀�*0��L?�\F�]�r^��"�[�_Nҹ��C��9�~��6t����#�|����i�Ȃ��Ih���AH�/�1�c�k#�n������6�C�f]��*�C`���S��bb!
~7��K�L�	g���1�;(ݙ�C4���ʥ��a��OU�^b�҉�����L׈���y��n�w��	՟�		a�7c3�� �K�I���}㼎Xc�C.�Σ,�mpx<�k��^���Iz����Pf�\]��0����\v��9����'e�э�]�U�C�f�p��(@�=!k��c�8�#I�X%�����X8��n�i��!h��C>{�Ye�?�׊4�� ���ߜѓ �(��`�|�x�o��R֍6��N����:�>@V�nr��$��!�{8�V�Ԙ����	9�:��)G��$xo����}�in����#/\�gt�Ԣ�Sx���������(�Њ��p3����<�&fG�.|;��ܛ#c�~U�TB7M���u1ȵH-���+����f�?Ai�Xe��f�����	��ƺ�8t����L{{?S���98�Fry]�N>rD�^[�Bп
^i��)^.�83��J_�T�(��t��5��U�la��fk��TG��r�W
%�������\�Y��糏qzF;��I	t�1�oiC���Ǹɢr4͆�n��t&-�yڹ'u? �m��dc��z�)ɡ[c��~N|�u>�����'&$HKҒP�H{�r	/�I^�x�( 'W��Ywj@VAo�tE0��p>�����8�߮n�h�\�P��t��>U�����;�@,��^`���t},����v�)����Sx�����'->d3����r!���6�~�˜٪E�RQ�њ�Q"�r�F�u]|�S��O��z!C�
� 2x���n:դ�[]��x��`ok(m2�N��G���e�r٨�u�_�m~����~��2�u��p7�ڙC%���sW�T)o�g�+?hpj��Ò�ȥ�}h���$��|�������*vCN��5�>���x,�np`l�=$� ]`B� ��󠊮��ڶ��!WFR+�4��y��q�	���jԌ��w.�Y�ۑ�t��\ă��>��f��������]O Y��(�,�+����e���Zk����2��\|���_���fW�s4���;*%��N:��ZE8�-��ߕ��z�Zz�:1_G�_Y<\`OA�F/�y�\�Qk��c��U�4��մ��t���� �M���6f4�<U.��dk<JK���ط��3�V	�V:�ae1Vr���dj����H$݋��d���v�Tav�G�h�ǌ���԰S�}�V��ar��y4��kHW�ǀ�!�)��F�6�8�;��]�~���R��yH��؟� G�*�hL@�$�l]�▲�%�IL��..$�# �rD���V�U	������ݠflS��Ͳ�P�X+���Te;�˩���d&񄡙a�W����_�0y����sK<������H�
����	�H��B<µ� �O���~㏐D��	YԜ"O�!JE8h�G@�}�׀U%b9(V�ˣ����,˃����9��h�*�!��jX�|���O���ᛕpʟ����}�7���ʢ�Ϲ
��{������[�H3���}�=[���|w�`��.E��G�]M^&�Es���&k�Q's-�0Er����0?r�ݧȮ��IQw�'��X3�Ů�*B��q̖�o��X:��A���g�*����.vJ$Yc\e�Ꟁ;;��_����q��_>D��c�L<�,�+��,��(�Ɓ��=�)*�8������X�j�9	v���Y��Ǧ�P�`�,ۇq��GN���	����ǽķN�Z�դ�O����[h�鵏� ,��D�y��j���|�QE���F��O�te7��Ğ�j2�7YTAgY�%�v��U�V-RG�����Uz��a#q��龴��G��/����rѫ�\�-6#���!����c�U��&����G�"ͤ>�X@�8��/��^68���l��}:�[�WJ��y�3�V���o��l�
���x�ygr.��E����A ճ����gW.��CA(��3yVN�闘�GU����Y�y�0��ժ5G8�g��})M��赤��.��=���� �->�c���K��n�ܒ�V�?,ԛA�[�@���\��S�޼��pg�·uj; ��73T�y����.<8e�vDN� -_��c�(E�s�}~�a�ː�J��-'�\HW���Hdō��;L�
�D��\�E4���8<E�͑{gS�;8ܡ�&�lEO��En��W���HQ-�4�ڶaΑ�9�l�ؖ�`�A��5_{|԰xp�t��� x	\h�� ���	ö 1Y=b&�D����on�]*5��w��ebM����{u�jQ6�{X�
��L$Ļ��ѧ���,;��><a@��ۆ�8��xB�(#5�H�K}.V�9!U*�P,�Na�J�l8ـv5��	��(�7�ǉ��0jt���ɷ��1� ���ǉ���Ǒ�7�{xA�m�w,^9�uHS!�~�l�<ɹ|7P�r[�7gJ&��x��&�n�7B�z'�/%����\�
�էI4j� 0��gO/v9���k��v�ð|�r���0)M���@�'���*t��B�Y���U@,u�Lᡋ��E/(��"��_;���]���8
��+���c�-�>m�k����w�P$��-��T0p�Gl�J�A�t�<s��vb7���C��f����5+���T#��}�?l�ŋ?찡����#LV|W������UҸrG�;>ϲ������G��_>bj�ǋ���*1�^HͿ�Fuct�Q�=�@i5�#����Жe�7�5E�� �0�1XJt�2��%��l�uv��K�0�x���Z ��}svӯ�2��O�S<'� ��,p��|��Y���[�E_@�mcFpy����@h6`r�1g`
8�	KV�T��O�@ҁ�Vs�=a'�>�.!��Z��:���︾�m/�6f��sos������E��aj����Q+8������$���͊��J���Dp�`_�`RH#��!Ljq��Oa6_���o?NC�����w^+w�����y�/�(-���<#<��W��^]�����)���eQa-%X����V�1�}�\��f�z]j�tI������ {�*�x�8����=�����$�+A���6�@����η ����H��!S����/�֤��p|�4U���A�x�Tr M���~��0< &1�����$��M��+�$5������t�CXZt��Y6t
_��Q
�],�I�ҦΓ��?o��%�R�N
<«�Ag�f�k3k��R�n���B���\��rK�jp�9p!�����3�N���̬U��ֳ/͈u������ z��h*�Y+���x�[��}�cR�`�-謰t��3�(~��F��Q��j��R��<�~�I�M�;v�>�Nc�e�vy�H�C/��Տ���P�]����필DW�Ժ2A������ӓYm��� ��18��I��,��[|�%���Ql��,�/�O'V�U�#�g_��B�<jґUh9�M��B �tvN�����:�.���Cs.��!l�~.:���`��*���Jpy��zNvc��Xx>|&��_��+ڃ�������ı˚�s��,m�g���rh�p�-?����]���BZ(2,����N	n��d���ʇ;�Q^ݵe��_25l)��p'��*��6��\c�`+���)�a2��&�� �C�Lh��\���A��� .�{;~��֩��rl�Ri�$�X��>]c�Ҽx�0�Z0�����������ٮ���=����� ��J%�� �=�9�9�Yb��8�!,���(�#9�ڲ��/5�h���L#!�!P'�B�:N�-�}����Y��a�b"_҉ҿ
){6IZLV�\N'�/ʙ�A�D�0R>�R̔i��4�tޜE
@�f �_ ���ͻ{�V�(��Gd���t��֨�m,T�J$����z��S̴.��tZ3y��h1An
+o�oae[L�!JuQ�4v����H+Fy:������?g:�9c�e�.)m}G��M��/��պ:g�VQ7;�U�fQ�<�CˬT��S��:*j��d����[M7�:l��S�tz�VmM� z��SA~_���$WV�h��KgVPV��t���q���K��e"�ȪYl\��s���0=�	Vm{�r� �λ7�¡�%���/7�Vq���]�py���<�3��e��FZ"�Z���)3�&&�<�	R��5�ji�2�7J�8�ـ��5�������|	�C�Y�;���Xd���#�J4���㐷���,���0�ۃ��8�q�#�8L�u��5P� ��FLJ�'ȩ�F	ԣʾ�A�`���á�y���O�T0~Б�ԤW���u�d75�Ш��;�K$� �9�3�0�n��/��AP�-�?���X hCȇ$��{Ĩ<��3oϟ�-��b�M��G���m��{6-,;��[��Nx�Aj��Tr�h���M�+$P�ԯ���
��� �	�ϯ�M�&���݄ �a��f���yPV���u��=v�GY�5���2y�c-��0��AT����I������	t-�E�Թ���Y�I�b�Et��oo�`�E���'K��g���n�f�r�\�W��\�ܟu��km�?8���2�������q!�a��!�KY�X����C]j� ���M����h'}�+eϢ����ai�~����f��F�/�v+Hy�����-l.�J�p��\s�M���P�AL����b�{�Ѿ��}��sH�,5�'5H�݌S������Gȭ��@��{\� OJ(_�2��ҳr_��0�Ĕ����;�g�u"�L�DI^%�������'�M���%:Z/�;��Z�|Ŧ�T;�.S�1�"N���I��GJC@^+Pz�OM���D�;��ʱ�U�e~lB�t͉���9-���������p��#�u݋h78/VO��.�������ڋt��=G����T���b'���##��A� �LIa9�Kɷqo������ !Gpґ�N��2�b����ZoL=�ʰ<��e>ƠT�6xN3[p���#\dC�@L�YL*e���s���� ��_�H0LڗS��F��ȍ[�=,"��g/�ǄC���C�9��rC�(
l1gpdѝW���Cw�̢9�Ȍ�<������jR�&�V˅u9{�9���uةF�e�����Uhgo@Z�����G0#�Gb04Q�ш�e�f����s[{K&�f�+���m�T�5g�����L��q;���0����O�o���	׺�nC���!���󻪡~"~���SZ��1��'��/&���?q} �<ޑ$ _a�1M��q��ܭT�_C�|w��!t�:��u��o�	K����J��'8��~_Y���b:'�&/V&���RZ�R�q���؛�e��!���4|R�졝��5��<�;2��+���{C��=�_u8��ɂT�����Z���1u��rN�0)�$�b��S�B������	*�R�yM�������ߥ��@y�2'�+�{q��6�����
@=�f�kơ����u拤��
P|�i9V��/�/e v%\V�*�����N�ܥ��;a4uZ;p���+��qw�K�_鉚GX�6wÓX�i DN����mA��=E{::Ir��!a�4����UD�uf����o�{��ĳ�wIJ*6�ۄw�����۶Y��,�í���b����Ņ����l����o@�[��
Iu]X�wv �sI�R!�}vN��y��K���K�}5��۹0]V��v������T��
#+f�p^`ld����KLq^���l˄�������N4zg1��u1y5�@���G����K����wP.�������Nz����Z�ku��}���_67�4�;e��,s$F���n�C6<	��z�Lp9�C>Z������W�}�&I_�5��>�׳>�.��_얮L$x-K�u�+�>��m#���{�{��4Oqd�nǴ���#A*`ı<�)�P3	"�.+����.��!����2Ek�Dgp�D�ό.�M�!x+|(3�S7Bu�,��YCj��xr9GK�NG"W@}H��Hv�Hv�2�˴�F �
lm��w=:������ҳ�K�_��ӻH�Y�Ɂp����x@�?H_��G������|�5>�"���k��s���pze.#��*��2!����iK�"(�v��2�ز��;��k+�u���X�`
�hHt����R7�k�����}l��Gԕ��,����}���w�,
�LAJ_���MNG��%���6*��s�
�.��ɖIg����Ҿ{�4�GTLFA{��d��[��;چ���2A�D�b�0��%Q���~�yz����iՒ6�ӥ�w�Y����4'SIZ��&�c�TK��} �X�6�o�~v��/z*��[)D[����O��#l���2Ց�6��;�Y�o�J௬d�2�u��H����KJU�4����ц���5�#�����t�?	�ߔk��%��?��*q���+�����!,f�B�)"�1�'��f'�s���
E����LA�}2u��9��e�_[��>5��z(Fv�t���O㟬R��`v�j��.��N�k����A�����Qs2�Rn�в�7����.��f,3����X����kB+�2c��s�C�)`��]ƨ^E�Y3Z�u�1��jɔ:�4K)-,��Ͱ��s��c -��DWew�@�bH�(1�VĕI��bq�T���#�i̓�Rp�o�}µ>��:zZ����R��!�M������� 3��]d�d��$�o�R��i㴺���DyL#��'7�f]׷��,�:���." e0���9%q�%u.���߫L���h�����¨���	<r��"g�H?�e����֖0�)i��i���
NS#~��jӻ�2b�čQ�?O3@�<���ċ>ڽq޺�Q�Q��H�$�%)���,np�I�Ǭ�w���T���� (����:�A��r���/`��8Q���|�D"����E�'6兩�y�S�[®�@�0�_� ������-?�z�G����$(M/�A��+�M Nv���^�����U�u%O�0r�ۚr����\?S���P��d�����PY��E�B=�(>�j�5-��HE�Y���6;�.~���� um ��7�O"��nz����8xE�<��C�Lqv����"^(M	��WA?4��3�;G�P����2_�������2�n�p�5n{<1�86�S^Y�<��B=slbuU8����gd����W�JiG��?����->�4W�<hE�o�
�1��t�E���b�E�Fz��� ���A"�U�OY��[�I�y6���X��`��?68�J���*!���&
>�/!e�QO1N��s�#�m1�,\	��؏�����)$�T�h���	:��9�C�26���"+��
�_T^7%c/�oD�># 4ig~n�Oy���}1�j�
���n��^��'��onM�����V\k安2b��$eo� DfeGG0$C<�p!�ѩ����#*��A�聽�jHZ+�D�3t��x�t������b^�4�SI���(����7�x�狠�w"̞���@���\ڶ����x�\L��N���y��͸�S�(��y����� $��9K�ٞE�V�[+�Za��/D'�H�1Eʷ~�hO4i���ͮD�=�ِ�A�|����z��;������#�Vꧺ�f�f�>��c>�{$M۝,�/���#���e���7��hݭP�捧$N��r�[�lb}"��9�gx��cȃ62�v����娥�V�M�Q�l�=,��C>�9�G������Vԁ��д+���nz�솆3��Sr:�nL��J���0)�����\STB��F�vjv	鐖��yD ]�	�]��:�L�}���Nę^;�z�\��5��^{�J�u�9.��E��1����T��;f#�x�hH;�eL��k�r�����<�mu��k֌�v�Nh3v��ʯ�zY�ki6�T�,a̖�窵ФW^�)���,�*����1[�Dـ2i�/�d�x� Fx�;`an�W���a�ԅ\y`�}<����r�Jܲ�Q��b��Ca�@$��$lm7?��^K��Х_�������9�7��+}����lhl������	������D�d J{O��9kAM���l�<�;�O����t˰kz�������Q�E�\z1e�R0�Z�2��`��9�^��F=���Zq -EQNݜ��*V(��_F1���Lr۫
K�&s]3zP�NnaL�<�\S�)F���J�'�Ѯ]�NІs�b!�9��{��E�1�����ɐ\l��x@W�Ί$�(.-����޲��<) ��eeb�ړ���ځ	�_��u@cE�r}Wh�t��T�[�(ه����:������)E��1'K�M/�LÃH�;��U77��:���*��/)!����͏�����
(�.r�z1B㰂���~M��ü[�zNh3!���n/~g`�x3��+2b�g��֢�X7�On���(��*>%~�ηf�"
gO�PBhH6A0<��h88�x��ߗ�hؼ�}����`�Ĳ��ԛ�S�,�v���'��(oܾn��U��������0W�!k\�eI'�7�qS�4Y�:獥�P�N���������h�JP2xb�QD�s��j�]����,�a@E�t� �v��~_k�.�С�}���Ԇ��A�����O:���KH0s��iJٗ 2���r�&���ȿ]��/���,o��O5xm,`'ϮeK����p���j>�H����!��\O����:	�+��rx7�Ee�w�ە�D��C���IK;G��
Ӑ	ڇ=,��(��2E2�~R���?��sc6Z	!�x^��YO�t���v�a��~Q�єH����!��8����h�q�^�wx%|_Q������6���&9������<�\J��Ʋ�t��	(OC�{�pD4[�_��wo����`=�D�"��~s�IkȂ!?���,EIJ����������wr阗j[l�~}�	FP���6��J.~��ΐ����0:'|!�N^���twM��ʌ
��@ ���DN�P.Ѳ̬�~ ���&��^�8�]u�`��JX;xB4�-շt�� n���E-�7Q�,�����iG��z��R;Q+��M<z�oκ�ԬD'N5�����`7�+ڦ���v	�b�u=\�s���+T�*Ρw���Kg��ePg�q�=u�@i_��f��܅7W[��&RwQ1�iL���;TM`�U��g�Tw�q���)�j��9�ωN����xJ;n���ܯ�G��^^�b>fHh�u��wLX̒����:r�.�姱��JƔ��KN7-��P�9�����,r�G����'��H�B����`f:�,�P<W����W��+����"���R�������ܽ3�/�`i�Ö���F��Q��@
r9"�X���@8p��Eb5j�����WV@�j��
�^{XV<�T�Z���\`z9��|H����x�f� �C��[+}�$����!`@�
ܗ��?+�.�*�/_�c���h-�ZJ텻N�{�����W=@S���MI��A�c�GE	��B�
"�6#"b�h�t��r�|���j$�E��$x��E�I��#8��`�$+�|�?�ȱ%�Jq�=Q?Ƶ���rI+����Zy���r�B��	���VS:L�c�^9�cQ�X�4�eÆ$z�E��X������8����+R>��{yӈ���G�U 0FG.L˴q�Zn`�9T`Pr���m� ½�j��wQk^�m�
N����+��)�f�g+}�0��Lmu�L�B��ƃ���E-ER���gN ��MU���9R)7-�K�[\�GlJy�HOf���r4G\:��S���{��=��0����^A>�wwL��K�0�s a��M����R(/�/ٲ�Ʌ���;6^�o�b���"r���/f~�?e�������R����
��S_M��?P���iu�8Kp�K�M;,#jL��H����m�Xf�`�"7��bY��az�}l�᡾�cS�1ΐ�bZ���t��>�$8�jN*T@ 
'F!�4�,�N��8\[��v�[.��*T>��IGk׽a ���X,�O�y��;���-tP��sa)��_�B�M{��&c�:g�����7Q�ؼ�n�����4I�Q����ྮH��q�}�,��y*GXˢ�<B��G��W�/sV����J�����6ݒ�$�ϐ��i7pԼ�A���X�:�۸�~G�0#tΗv#2�3��>ES�8{�cV΢{?	d�[K�5�q����ݭ�<��]Sq����\;r^Q]}��rD�b���W�ܫ�*դ���z#J�S%+-g���[\��r�I�،T*�r\]�=Sb��}�%�o�w
��n�i&��QJ耏Z��=C'E޲�A�АS�wH� ��3)΃�M�Ls��&�+�5I�Jt��1���6?�W��o�Uv�_j�ӚTӦ���ض8�c�_a��B5�̪��Q����%�FqT	̏a5Z��F��Ǚ��y5����Q��#��e�;�.�X����/T�
���G�w&hs^_x\<5�q�3u��nAE(������p�*���E z�v����=[���wq���d�f��ٸ�,c�U1�Ihv����lo�c��C��^�O7��oi��l�'� ������t��!�����gĢ
ߤ�)��f������qB��|R�N�ڝ����Y��{���50�YK�u��EW���DF;���N�˿h��m5K�)DS������MD��!�@�����&��4��,[��/9Ǫ��fAʆ��z��R���寇�
µ��(���6	�V�F��ɐ����7�k]�4�� ���ʑ�d̋j@���bR/�V�zL��i�����zN�NR�9c�_��jJ���S�Zq��ԗ�n���5�daqb�]����N�N��*}Q(��;O[�^/Z)��h���,���;]��S������m��k�y�`Dp":ǴC�|����dDB讘��#!��cZ>%Z�J0):�mT6���"k�,6�vP������w���l�=jw��tўVv�U�-I��-|94#�9�?b�\Ӭ������I(*������֝S5���M���1�}6���"csG�h��^
��o����ݵ6 =M��L�6꺋��j��2�6��Y��d����SP������SR�� \��jN�#�����H��Cw�Q��.�RN��Q��z���/��Dք��p�3�R���gEq�z����
K�������ap3���=	�/�&�m�q��]ʇ�,����hk�J�գ�/K��N�fC\����Ab��>���WQ�&6=:׷7O��/p�e���B�N��u��Y+-��i���o��,e���+�7L�s�%���M���Ɔ�]�6������߫��δ Y��ӵϹ4qd#6��K8�8��l�1�:�稆f������
�'rծI�1���2���#�l�\a���6�8�o��ѿ2X �1��'�9���m&a�W�����i�0�����;l�xP2V���g-����!W�\:�wT���d���+�I��1|	QK����r�a0��x5nۡC_Jo�ɻj�m���F�BÔ�Wa�E{ީ~١ׇQ,�q�"�>Hkj���fU +������u]�_�H�Z>����bMD�{RS֦A��a<�w�++��V�ӱ�K& y�U|���t<͡��.���p��&-�����T�@V�s���_u�_�;���+'�~y����3�l�iy"I/7���r��n������8i�13���'�%m�e|����M}*�����B=�{G�x�{��\äv�_7Q�	��H0e7Bf�����;h�x�|V)f���b闥�	4�o=� ��m	�	]'��6<�rM�|OP��
�%����Dq��,��6��4X�5�C��I������3/�<�9C �~v��z�wH��y�|.2�������,g����fA_B�����f��ф^����Y�p�ɼ�q�V']�@p���/���wr��	ʺk�U���q=m�)�i��o���[�j��4�CP^v�p�$:�-Z"��<L�>V2"uar��q�H�{�$£Z�	��3%������D�s�ƿT����z��,�JBI���}�*G1T�I*tcF"�ø�*��^Y�Q��ݞҭ=��p&[>��SpJ����$������P��K�wo�}�OS�{B+��B�]��]a1��J˜l�v��Mg����gFkt�2Z<��NB�����F��RKU�(J��b_D�_�-�X�ń�E&,y52�Ż�	>��S�LǇ�Aܟ8����͋;���z��Jz�Y/��h-���5Xc��a4*G!P��^�, z�+�]��u��D)^:;}aoc*u@�q2�2b{��E�H����%�L�l}�f"�@r�~����uGSK�&�l`w;\��_��M�?�ưj�^�~�R[B�բ�ۉɏ��r���_��PAC�J���[y-yN�)W߻��dN�����퐮(�j��������N_�l+��Y�����͜���s��O����
�a�i��x��vVQq���9�z���X� ¤�γ=�ZdS|T��g�9P_�+�<�	NP�|���`�[�	��ʴ��F?���T�5��|�ӽ����B�z�O�m�3��������pdk����Nr��{�cfZ���3&��C�= n�?���st�sx��m�� 0��b�Ư4Ӎlʹ^�ɮe�y-b�
�T�ҶP�Pq��i[F~�Ѣ$K������ö�S���Zl�=Y��r��ui��乏'�Y������kZWT�';��a��9
X SY:�家��7�(~$��c B����	O�����!��vv3z@��?�q'��קsГ��Q��D�,���]�!ex ��ކ���֚Y�x���J#��c�ڀ.'T����)&J��	��tr�]��/�ܔ~d���ہJ�D��6��k��)���W��������J��ǖ��=dG(\�9ҝ��m���4:������2�(��HUu���:��6���5�EP9gSz\�kR<�)�=I/�uſ{��jj;�H��0��$5��"��<#�����^�7�9��[]��*��"]o���2-3KA�t#��V�O��l	�y�_a.�ތ߇y6.C�ɾE��9̇\gN��3Ǔ����
������U>�b�?�D|-=:���.)�
����_@=z?�\Y��̃�"݆��X:�b�ǃ�!:��FO:�i�l��L���P>s�`KԬz =���@�>����L��x���-�E{�k��ن^1�&���Ƃ���Lڣ0�#~W���İ��6�y�~��^[K�{N"~rd��m��Lۨ7%{�)ȉ]���న�P��7��D��gA�(ź�?�� :�8�W3�O�D���&���o^����Q�����v��]�N;����%i�M_���q�hBa'�sy��\�!k����+��x	yrz�^�K7}-F ������*E�� r�dDx�?�i�Bډ��UtW��q�i�����Iݲ⢄.��s1�M[X�I)�ޠ�BBԻ�0M�O��������l��8�E��3/����Z�=�+�ʳvUzKX��e�� ��Th<��fƃ3D�d��1�Ϊ)�ufDr�G�JvH/��C?.�M�k�P���I����݅�*�RnI��m��[c�ܩ���Z4Ћt�G��0#���CҒ�ϩ3���p]������Xyz]<A�!j|5�d!B��}�Ǭ<EU�tl���_�q�}<��=t;e|�C�g�:��{��m9�L*��[b=�3�.lgݓ)�o�����n6��@r��]������p���7��'���o�~H�Yd�m7'�[�q�d_7�F��Ph�/%m�
ԏ������g[�э[5�df�y�~�̳�"UO���V~A�m�̝�P���@����Z)2��ő� ����T�����ѻA�	ơ��K��G(��B6p��7�U*�8.}�ֵy.���qEzn:/,Sb��G�!\��T�k�Y��.�^���P��i�v��P
�9�IaH��o� �4=�x4��\���6)��K�:[eri��E�?x��4�t~KQe;�xPc9K����I�L�_���fJ�9ςP�RO��������/���g̡�{����e�׌vYf�*��o<�����|�����}P[�� 2�����%�Ez�n���_5r�28�O70�ȿ���	�W	f����X/��nښjocܑVnY�N����q{��u��F�����)�G���Nꃴ��-z�H>:z��;�G�e��_
��ub$��P�5Ւ����-��(0/f&]�Z ��m��.��U�{|�I��r�jE��17o�U�2�m�dF���G=8v-�W�<�ΰ,q���$����wۖ��� =���z옢��یemƟ��A�ύ��Y�^^� ����j*!���u�fԦs�_�a�]=�8sF��9sJ]�а��b��5mV ��`��"��h���\�;�Su�=s�w>�r�S��U��м���e��� ��s}� -���x����{ǡ�C�5���L`	�+�;���XM�W��h܅��-<ԃlg������}���վ�
:`!S�}�e�qgY�B��{$��B��'�p@�6q�f"Q�����c��"f��L�C�>�atu��s��c�9�cU��7�U%��oh����]-�=,;ny�5jR孠ݵ#����ZϹd WhS��P0[`���~�+��Ž�#y=�y%��w��H��XrǗ��g��7��9I����,�$Ŋ>����K=��ׂͩ�s�颈~��A��,�}��]9l��'�N���2�Y�\햃�=��J���[�>��a�%&
��V2���]���9�̝I,S-�2
B�{?���#���F`�i��W�}#��֥)U�`���l�ܲ4v�������ףF�z����z@�عD��B��q����ˍ�Q�)�}��ho�h���[��u�HQN����j],$��(�_�:J1֢��fI:�»�<APZC(�w
�ݰ���������/�u:����2�W��7.W�̫L�´,^_����XMf�L��^o{�ᗓ;yˬT!Q#��%+�	���66p0�5
 ��i+5!�"P���]��9���š����Ά!��8]X�b6&�
��6�$�2�O�I,�֓�I���{���#ime��wYG�zά��0x�0�T�j�����E~	�Y�*���f���؅��g ���G�3$~[�::D9�h���TM2Z5-�ho��N8���-(�iss��f ��GtldW�'|�o=w�:˖t��L3��aՑ��}�b�h�^b�h�T���8�
;���Mxj��3̞i\F����DN1����:���Z��
�u�aз�_s�����τ~h��������r� %f1�,�i.�T������z�����:��w�����e;L��g�d���n�`¶;Z!>��{v�MU���a�4|��B@Q��ÇQ��׆�N�)�Fb�֒5#vj�
���c��U;)o�3�5�2U�&B���)��c������b4�X�co� �Ej�(|,�5*����>}�f.��UhrUsD�� ���D�d�ԸH��ր�"����͏�IA7Ӈ��z���5�v����}p�at& n�9
�݊����6�o���T�l�K��`-���f������}
��w<%S�j?]��
5�3Ӽ�͞�Էb0�V��Tg���گ�lc ��4�@�C:��p����
�l��e`0�=�8%	6���`�s�+���Q:~zY�R��,N��"�	�2�� ��Ҕl�>(���`����r*d����7�z(��RD���ֽ������`�������ka��s���f���/�a��c��oN���G^�S)�W�=�)��e�1N�0����a��'g�z���~q��RV(j8�J���z�d�)�]�;��9u<M]@�^F���q"E�4F�Q\54O;y���l�͙���
0
�a#��x��m@Pz����$�3����}W�?R����xf�ǨL*�},AX��7ûӼ����;]M�r��c#s�����(��Y�Kcd��[�㽺'�M�g]�@O�%�����C���5l2�7-2e�}�R��k4�hdS���cB>�)���@���t,�8�l�ܾ�(�B;�c��/��5����hre�sy�fu9ؾ>a���<�Y����{.��.쨷7�u�O�Ǝ°~H���6h�.�s�)�e>A�F[��O����]������T�M�y�[BW���?��|%7�'�X�������{5�RZ��Q$3�*Z�VD$î�p�_���A��1��_tq���B�iSĝ�.~�c'��y�4G$�	9j̖�2�Ɏ�t���$	��>5�
�:�pX(�vŹ�]���j��v�/��s�����}�Q��r@�φ#m��(;ED$�B�ԕ8������G�ˡL2�H����H:#�Q
�W�3�r1ΕX�>:�	|��~��j�Q���ԓ4$)ʕ�{��G�5�'ڸ�;B2ǧP&.[�v�u�T��֙V�%Q����C��SJJ����xF�}�y#b#y�O�׳�^�1�"/i�"����+U�NC\Y
����w����!H�%d3r5>�[(�;N/�OTc 4�T�;"z��^���W��\�g~b��"�8��Z��7��� 旓�\{#�p6�O�����L�^�z�8�@�e��N��3��A��J�EDm�MG�~a�)7�a�M�s�e�| ��DْiҴ+L�O�93"�� w}��� � _�a=��-iv
7�`�nm6�S���wF7Ɯw��q��=���ԏB�m�T;mS�<��U��\�V=� �SH�_ŦvE�.�_��F53��]�5�DDVl�� �|�qM�tү+�M�w� |�*g��H�6`i� xZ:�K!�m8LD#m_N.�����<��q��]�D�2�C���t�nV���ζB��Y�G��i�ҙ�hx�1��l���́K�v6�QXA�"_B�mAC*�+ ��%b		���x�l��oj�c�	|CۥGQ�����͟��2���ҩ*ӎ)0VS�ŉ�'�z8�y��nu`�iANOr�����kv�*��a�D����k�j����&�҇.��oFZ����]F���]��gR��^����j�%B��� �����R�@��$<{߶��^�'nfc��ƺ!c Sx|p�PӦ�D�ed�A��>�Զ�)�U��u{�;��$ݵ:���l�j��p��ǉ�Юa���Xbqv�%�TrDf�s���7?�	�=jc�����g�ޡD@7v"��S!�y��f~�(g��!\���:m$0g��ףs[\�Z&���w^������Y�`1�'�1N�������l����U^C�Sp�oNj'�PD��j�=�����Bn�Ont.���Z��)*Ӽ/���R14��ըPs�l�DK��)���%M ���,"�E7��x&F)~�fe��@�����7�z�aԻ�G]���1?&���I+�PG
w��d���ˀW��tלx�t��L��!Dt�gԕ":�%)y�����ʵ��r�� 7:I��-��@.<s�s�_��|dQ2�>er�V�J��ދ1
�s���A0�P1u��y�S^�?�̔�'n����rEz����	���s������E2���_3��3�G�͌S�2��{���)�L.��/vb�nO1�L_}����(Q�[�
sl�{8H|�臮C��P��E~eK�R��h�{&��9�[u���6[9'����"�y�~zaX���8�:�s�֏%��I�8�ê���"#~��q1�� rN�W��G�M��-}+����P�
�i��_T��A���Թ�_��Fꨒ;߻��E��^��X5���L�$0�\�<UM<o�W�/J��Ou���jP��D�0�V�*�g����92���H����ل.���m�es��y������'Bm�b�!2�BԸ��)�ގN��mCG�9���,�/PG7)}�O�'�l"�wZy��Vi
{dx ]]�
����[d��@!�6��AF�z��X�'g�j�����,�#�����.���L�4����7��=j������Y���\r]�#H�����.�_.mԜy׬:��o=rB�
:/a�܄���I��
B�ɀ��(%�B�'�^��9c]?eMq���M��L�ܶ�F|D8�����\dT{`��,�ʝk2��3�H	�
b �fv�jz��b�,�t�)T ,�9�Q�2	��BP1��_�oW�u�J3���[+���W8���X׀RZsL��J���NǼ 4v����`����D����W����cr3I�|lk>���ϑ1h��C��wζs�j��T��Fu�koC�`p	c�hNj���G�����Em���*%sK��)�����m��c�V������$�����\?��7(g ���6�K�<D��EO1v�_e��lǇ��H{K�<q�ڇ��@]V��X���j��ZRp��(*�l8��Ŵ.�ZBV����e�\m0�)���1��D�SP߻#	���<���V����j�n��dz	G�����6�+�˰�_�(٦�l,F�5�B��aC"�A�L���A�3H�,�.��$B��Q�q&�-�-�JS���2�x:�q��2	�c�f��s�1/�ꕾ,Ћ��@�/�"Ϣ�z� >�L}5i?� Vw��7�5 �"��e����0�q~K�RL�	$𚮍}j�\)��7���r���s���56��<`��Mܗ���V=�rhw ���z���^A��[W�`f��C#L��w��(zyT��.PƹHf�� 8#�������Ɛ�Ȍ���m�c�2���ɚ;��K�5�o��}��a�񖐵�fs�;9���"�Мف��Bi(�G��+|��"u�����E�����Y�Y_�sYy����9��z
c��oj껺ƭ>aG�a�$��� =A&����r8W,��9#cU	0.��>�����텈������������3����ƪ��O���A�0��7�I��0����p�u���>T�tRg��MS����VB$�T~��t�)~�v_1���$��T)ܥ���~J�-�k���:Q]�C*b^�&�����x�]&�:R�Lה����C��\��W�P�~|��r�m�uH�{���j��Ey,m����.
�y,�:_�e@���� �^T��z�.�$�r~�%/����@t���K�u+W�8�R��򟢯WF����1���R+I���!4��	Ă�۩ջ`Q��⢛�]�	z<��/���{�e7����e�a�e�&��wV_����Ձ�cP�ݗI5
+��w���g8�BM4�^.`��:`Xh� �P\tD�YA�j���I6�{	K��u��j���.AN��{䔼.)�#��NڜN�.ax	�{g�,��π=��T����@�7����w�H��<�H�i��,a���ۅ�j!�3�G)��g	�3��u.���)�Y��-h�U���ϓ�j܂ª�(�HQ���ΪMcj İ7���W��/�72{�[��8th=Sĵ߼�Qn��E� �T'�jQ�.�i����{(dJ��>3�ӫ�8���hR�K��_�Z�i.����/�6��}9���8���c�8g����������r���K�g�F���9 6��N[&v��'�$��À�j�ʪ�|�=����Q�͕2F
�Vh�I�����Iǘ7�̉^�v�&�z��ZG�����p෦�u3mL�-t1�ף��m�ܲ?I�ʺ��.��>V�$�Q>�^�M}��[�&�)_
�+w�(�'��y^�@݊�횫#�����>�:A���4+莎t\����)M@a1���N(�ޓ��e-�ܲC-��֚[�%�NƖ�}����a�2��g�?�H�z�ԯm��\z*��m�o}I��$� �,�-@a!ER��m -�c1�(e�L��u,=�~<����v|�;���ȣ]:�{_�� \}ɱ��r������u�/��U��sP�:�\���퐍�D]F�v�U�?��UQ7˽T���Ҫ	���|���瑝�o��,#��;��N���Rt��1y��(��g��z�\����[��-C-~�-;��Z-���l��R#���{�v�9���SZ��^�񐴿Ȱ6 �a�0;�fl|�U��(B�n�C,_"��D�e�X�`C���&)(���o�����^��f��5��=7<�1W�(�%�	��$��-.N�����3E��Q=}��yQ��B�*p�g$ۗw+��dޕ�>+�+)�H�L�h��b֓�n��s֠oV��ڷM#X?������2�S�*P�0a(ٗ'�l5�O,6���ʷ*	rB��X�2��ɛT��Hq����c�A�Z��g�r)��>�i�����u�~&����y{�a�LJ�kP��~
XB8��P�տ�
��C*�.&����.���%�}�e��M݇"�8<E�����kO����b��eT�����ѓ�g^�4V�R��xB��d���fԌ��$���n�x���z����)����3��wL� 55롴`��tr�Q����'�[��-X/��N���[-I�h_6���u�X-�����=�&��j�j7�ۯ1�~��-��X��xّC��|��[ٹѴ��`��_R�y%�:I���{ � *{��bT�)�K��h"$�95���}��k쟉� ���;']���^�/��]���Wٜc!�����ﯙ�]��|�^�4����h��$-,(v3��.�'�n�Rb{`�C�Ota�����D�p���r8eڇ����X��'�i�!92�
:���*M0R��������D��e�Ozl��݄Y�q�#y�ҭm+��ڳ��Is8����s�. ]�B秥ٲ��YNk�Qw	�jH��ah�`|�yt ��[3$�{����l�B<����p~��a�^��\�J㟆�^D�d�G{إ�j�&�U��<z�P�(k~;v�4��u5�#
x��o�?Ʒ�x�K��:���S�0d�rQ�$5���7q�Q���Z�e�%�P���.��r'���~�w!�i�5�����*xvMx����yys��A�];ض���\59�ЕK�\&��4|m��ZA��,�:ｕ��Y�څ���9w�(�P"���1�gķ�t,�}@gX�쵲�;�;��ޚ��9^}���m���������)��3XГ0��p��s	$�ݶiB���qm�$�+p���8G�M3!�cS/1�����@���p��㊒p�Q���̓gL�|�܅�A�2��\S��r>#���z�|����ܜ	�`,{��L"�D�H"1Ԭr�#�゛��� H[��@-���z�ٌ<��>�a[���)x���*��,�� F������+rNsL_�b�{�5
����*�����U@(��H˭2��l\�Ȍ�d�Zb��)ϊ���+������6�e��	.V�d����P���Kn��d���?�'�6��)<�s�t��@[�'�W2=,�A��4�lچ�$�:O��G!g]����z��6`�|�������X���l��=J��8�j9����L�'�S�������m����ϯT��֗3�/���J�x�;��<���\q@�D�;����N�����?/t~�˅K�<x�
�pIn�`��a��!�n@��cKQ���*@���S	��,E���^9@˱�W��co��Θ �wR:����#c5�|���[RW�:�N3�%���Y����C7��i�����:<ݑo�# �rM���)o�>�X����(Y�����K��P��m���4��=�<��{N��;�P~�{���x���i���}��_h{^ptw(��cx�R1�Eё4��Znk��T�����]h��s�I@TRS�%$j�^�ֆ/Q�N�,6���A�\���Z1W`�׽�s��LdLY+�ݼ�B��z��c�C;�Gu�Me�c��odR)ٱŉ"�e�
�J���^�!S���ls��Ԙ��S�����������r1껕!^�����O:�����j��a�C��3��faMd�F���]5�X/y�nɣ��e�'bw?]��4�=3h�,�v9��Z��=�j���||�^�P�>��B�+:e�b�B��@�*��8���pϬ M~4����Ƕ(s[�ޤ�	z�0�t���?�g(K݊��b;�����-�y�����*$:,���������o��7-g�L8@�$/@�t��k�~�l�&�o��߀?�D-YT�m�3�}��)�`�M�j�e��3&�K%��I�m9o�ҽjVX@j��O�;l�������s]���t���Ft���Ai�OM �b?����˫��OO`Av�0}�^���^!���D�8*�>)F�y��vy�0��c<�0ou��1�N�.�L[��f5\s~��%�ڐDK���#����*L�X��۩�Zh��0��ORt~c��	Y���jXШ6�+걺9}b2��s��~�lr���յY�ׂG�o=[ӒtYps�(��!�EMp����FC�\5���}�4\R42B��i���h� ��Eg��߶�q�D�{�_l~�"�)xǆjRb>��h� ��rd2A�C�%k�Z��_�n
�l�� 
�{����Nd�)�(�Ҳ����G�*9M���YhJt���N*���^�jpbL>;�1)�R��mxS�0~h[�ī�4H۷�I��.Ԗ����2.���?��"���܇����E4[������`��	�`Q�L�`�4A���?���nj�6������S�N�W�yu��<t���(�c��PЗޞn��GC=Y�U�,z�ʊ=U� �7��%ZL�F�M����ɉ�p�A^�a=���S�%����%������}4�AC���*�s��^݋�2.�骲�VH�u��ɞ��W����7?�W���>ۼ��	��ԥ���fƨ�~�Y~+��<��H�<s+�������l��%Y�17
Y4j1�Dwx�u��Л�_�L�8����Y���×���o+Q	� ��3�O�%����J覽R��-*HQǪY�r���|�Z�!g�v�D�w3m�w���2�a���Q�[Fbw����o���K���5"i��� T���<�s	�Ax�iF�Gl#���1�z�b[�@`����G�;-�n�p2�{�,�A�;�T�M	�/]�P������쎲rK�pm��(0O��IA"f�Wd
ٞ;�W�g��l���5� ���`��
�>�!m(�=H�6�������I���1�T�P� ��3���c����Af�[�!�?���R���y@�(��۰�p5g��U@-������>�x����LAE��0g�a+b%�N��h��F<���w��d�Ƥ�����9c)�BF|�;��u&��;]q�Li�Y����p��Y����2���Xq��$���׃��2k��l�%�
�Q�.�;��ro˹���<`����y���:�g���qc�����5?Y5poPJ@�	x���͖��vB$������{K���%N��d��1�B�B�laH�^�.�F��M��ҥ�˟KM�}N*�|�
  �k��;�c��x�����߅�&M��g$��k�,���&c��*/z{�Ζ%οoM���V���/z:ht*+�mr0#���;���U>E&��ke05��Ü�ff��G��Qn���A�g����9�V��Qv/�[֍�e�4l���\s�_m;������d+#q���sg�Q* ��\m�7�q�V����p�|�5��7��E�Գ�@�8���Y[����%.F!o��I[=�� ܀P�2��|���	�p�O��R�(Zw�[r��e�N΁�	�$�hH�n@Q3��P+�_��������7���8_�e�^�!fɘa��m�NqW�������C����P���s����<n��O�Z_B�8�G�������"Ÿy֩���:�!R�G�̶�ׇ�;�3���\A.��@,�����V�x�
���υiګ���e��MM���<�In1�TM��9�Vz�O��7.��cZ�]˲$nC�����[>��"���J�u�T��:-�Ӌ	<D�"O����|/ig.�zF
�G�r>+�BF�5zk�r�;��ڙ��#� �	5�zۧX�2���=��-��?P��Dϙ����������
�G��y����z�G_�;����jM���W�E�<�Ɗ�ՀP�ڵ���z[��6�G-w?l<��p��-�����w6 ?�>+��m��;r� ��@c�8osQQ{OR��W������VK��D�8�oF��z�D���5۷���ˬ?�Ub"`�Y�-I s[��<����j�(�f�-Y�#*%�Q:K'�q�
���y�_�pa;�/���N9��@�<ƴ�@�9U&��o�BӠ1D�N�;�$3�U�k�(��z�O��+�琻5=um�c΅ߘ%��"�B*���`aipi%���)dl�=Ħ���|���8�Y�@���{���szL��
RJ���]:t�M:C��f�5�l.F!@W�"���Z�4��c��ϓ�AZ���@fIc��.��ݭ��G�^?�d���ܾ_gK[`]���xH~4=�+��<���o�Äp�>*��Ⱁ RIt@��nsܔ'�7�v�P�����/��;�G�fq�K�G���Z��Yj&_+�/�����L.�5�=Bn���w�_u�qV��0�>�el�Q�2O`��jv@�tH��E�V$�D�f<1�jK%x021t�S�r��6�¼	 "�&~i�m�|��k�WI�©��ss�v�
z�53~b�Ѷ�*#l z����
�iT�� '
�~C}����kĚ)i+�E8�5Ve���y���Kb���YS�}x���/��M`��i�9��E��^t���m!S۟��� � �#�l�������x��{0/V������O_L��t�E!5
B�{��	爁>4,;��rATmV��$b9L=�0;4/�-\C�U1LE3\���y�?4:L�@����d}���|j���%�����1������p�z�r�i�(Lbn��8�����1Mz���63ӡ$_���h�>�����ی��Ui\��p;�y٭���g���⇏v)E�c4CD]L���=��9��ua�F*���2���U�f��k�hV��R����^�7`���3������jb,�v^ذHz���ϥ���b����X��6n�p1R���B#�t�Fw�~�4�f/d������&�'(�W�����Y��}zص��x�vk,P=2G�7����'��7˙�<���|y#��mw���Y.�OL��w�	R�J�q�)�*G�DF�i�.�������	�"���+p��Yt�,1*�	)�q~{��*Y�;���M����Ow���;o/:� ���������EA���m�z�QxɌ���-���_?����uxwؤ`�A.�	X|���R~���@7?d"�t�U����C$�����^�����&���u+��G��F?*�f����R���S�ڥ�L���l����ILqy���[>*E׼���M-�cP۴xY眧-8/j�ڽ����r��"LD���E�1�]Ӛ�\ mD?����kP��,*vWc2�d��0Ӷ"����G��P�����T�k[����{����� ���+&Hl��dl؃���d��P!Skimo�dl�s:���w]�Pmyg�IcG��+�J�:֘�~��`Ԣ�oJ��y<��Z�NƋ����s�Xm�z���&K�K�Ph�-4�q���~p��F�������!jj��V:-�@���>�<��R�E�!\!]��ִ��ݚ��#Zn�qcӛ�uZ�iuE	W��eƌ��Uq�A2��c��5�1���z����A!��o�]$q�<� �s��v��{a�m,,�>Z�I-��>�29��0�h�be�����ǦҞ1�p�]G�4��[�vz��Y���U�;WB)0�shj,�i���:$$��)w����R7K�n���<y�۔�\�'e(��|PLG��;;V��D��,�+D���G|��f5#m��|˟Տ�]�|�zs띳8��~̌�#VJ,DDDa�v�Ȉ@z����0�
�!7�J{72��}�T�-�����feeŁ�bNW�HO, �4(G��7� ���vA���i������O�0ZG����!���ښ�� ���������\��s�8���|��ۧoǗ .��5�akC4D�%F���`~R؄dx�U�eqJOg>����t�N8'����T�dK���_N�z�]�#}w��6QD*���Z��W��[����N]0�߸.l �S%����H�g���`b��1$����?	/S�j���b�oS��+�~1�h��c=��q�e���v�ؙ@��i�c,������I�x	� ��LYfϣ��4�y��<VN�o�P�y{�on�+�D���NԄ=WC�F ����O��Ev{*A��K�҉��]�HClm�\mB�fUiϔXx5���z@�Q}ڹ!̉�?c�l{VeK">��ƣp�p�#Gk�k6�����^D�_�$v�"���}�G�+�Iw�� ʲy�E��4�҃�i t�	E١0mRM/�A�������,�e(�����QR `Y�0�h"����D�r�3}Ν+��)|6m6�f�|�D�x�(�^�
)e|q��Q�\��7�^�E+a��q�Oc��!���e
�Y'�|OϪ��$���t�Ni�:)��a�	W_�LS/ֵ�6yI	d;�D��
jC�>�N�a��V����-���{���bm�����"ӓ%�_p�p��E��4�=��'4-�sѫ]������]X�;C�gۨ�i�q�k� ���ڔ�2�S5p�V:g9�X�	4]�kY�y��D��J槎<$��^xt�l�� �T���X�@Y��G_�.�Ζ��9�SGͯv�W8�ϸ49 |4-*A�F��<d1(b����2F(c\9�a����$����P8��꙳�ج����O��T�����|�%Ҭ���۳�scK��(iRI{W��c�� �IymrU���su�f�C�\+�vQo ����?���Q��zc6eO�]�;��i�Ź%��z$�%�)+[¡�?�gqq3�Å�b)[�Yұ���Kt���;L�,���@,7<ġ&?��`���)��#��eF�AA�Yŕ�u��w�� f��#�o�q8}Na�� �z"�ܢ[g��ㆇy!�'я�o4)�3���cӔ��$ͦ���M��>a] �����7���g�]���h,U2�vDؾEHT��Y?�[�o;���Y��k�S��B���'c9��+ ^`R?E�U��w�7t=��J�ܖ���\�Ld���%�Y��kɮl�/M=�h����gw@�Q��<i%wu�l�����z�O6_¬�Cd���%�����ysU1瓑HK%��2+��𗶜S�jgG�'�{��ױ#�Ғ���uᝂ� A�`�䣬�&L*�0�x)g-�O�Q�5sf�D������?��
yf9X{F 9_�8��Ɲ������{� ��p�0�)5��[dU�����ģ0Ă�˵�l��f��ˡ6bڤ�7$�+�aY�:(u�o��n�.��/|n��V+~9-��̖��ge�]�_�!_���̯�|�ś<�a@���g��T�Ǵ�@"Z��/�)�hO!�Wė���qsg�N�����}�`D�=F%��q��u��m�UW4<95�5��j��Q5����W��$`���u�o�/��B$��ӷC�_��X-5���.U��_oh�71�0����[�/���]n�A�_JȲ\;&�c�2@�q��V/���b��IoR�i�v+����:�l�u�.����]x�Rû��?H(�[��fV��Y޺gwI�u���Y ���_�,܇@Ӫ�F���rW�Ā��B�>�P�:z���i��T�BQA�V��W�{���1��2�e�@*��QoB�N$�;K��TLw��j�N�B��N�G8�D�����Yw���K,��1��m��)�����`5�'OJ�T ͊�s�ÿ�T�f�ǜ./])���Kn��F�S��A�! �C��)���+�{�7}k�H�ɼ�4��1Ia�B�P�ա���D��_���tW��&�屃��UN���:��F\Lj�_-w~V��s�{�h�``>>C���,� 녔�v ȼ/�a����C�
ǃ'��kv��V�̧���}��:����n�� �lC���@��CeBJIzMv�Q��ld[R�����4%�X����Z���<Րd[�:!/��qL����p�C�I��#���Nݗ��U���G�<��)�3�Ӷ������"ݛC�l�1��q��]is��B����
��c檈R��'��=���y������~kc=<��k�8�����I�J[��Q�,������i ��p��e�So�ZM�q,.x� S������R�v����-�Ú@��oU��yqkŃ�!���j�=vAzDwvev2�SQ��:lHw9"�����p vD�TF^ߒJŌ���N4w�g§~�וM*Y�G�Ɋ+�c6����������ю}��`�t���(��xB�Zc��`�c��L�;�CT��&Y��KI>	��i�8�a���Ф�fUA�$$��U�fb���NW	!\'�,�/����Z�s'��a�j�����Q�M��!�Kԑ1�q�-'oPV����RO�j�@���o�sG�8�}��{�']��\�ڰ.(?���F��^��������m�Y�[�S�:%ż�����{�=D�*�eL�`�����4l���V:�ib�W�yb�wZڏ�u|x�F�ei�D�se9ϼ�\�nk��Cs�?�<�h�Cz�� ��@��Yۨ3k��|o�x^%O���Mبx�g �;�=�4��2�|�?�L�:q;eX�i؋zH��q'���w�����O���p�,�N{rſeG�M/���'޺?�6ު($~p��*~@٦����<��,H
ڬ,�&M���+׈ XT%��?BCO��(���b���g���"T���K1C/l	��{?�g\/�ￋ�eP����x�_|�P%�e�mL�(̾7�@��Y�|Z�^������O5Y^GW�[�<Su�c����=���4��L�2�i�蔢�g��w!�n]I�k,��ּȯAHz)z�����3�4��R>�+}�s��w��a_��Yu�}������f3����i7'����L�#�ԙɰ�Q7X���7W,���@�/��~�����6E@O�1�#��I. t��V"j����fR��1���QЋ3x�B�����G0==��z�UX�n�?,���^o���eW��m������-1O��E�v�E�耊W|�Y'N�9��,~oq�gV�n��Ym�]z�7x��H���C�4���9�z�P�<�'�u��j�a>P���|��rql܍X�̘��^C�����o�Eo�r��ȓM�-{�_����
Vm�@���o]�pf�sZ�Cp��f�F�utx��B:mЮ*�o�iu���rW��?k���=p�ݒ�ׂV"�U7�®�p�/&玸�P���?|,��5�c���k_sRUɖ����)'l̜U���Z����m�I+�Vx�6}�Q492�w?�\����xѻ��l�_�	�	g�f�B)��UQ�qEiQ�l�cR���3O:⣲��\&�i0��� ��[L�m�L��'4B?f��f�w:?|� -�fc��΍�: �5�l��� ����$g�D�u��.<W�8}�J�ȺP��٥W��<x�B�g���]$�����"G�3�p�f� N�_�|�PgkO��!���{z"҄g���:��·�jc�?�� �,ˋ�_�}|~Qsuq��u(����5�EueZ;i��Ǻ^|�y�rm�i���0��+�>��������u�M���"|+Ap�w6� ����4snW�j�?�b��^)���}�[�EC	��hk�%n�8��Cb��x_�p�
�A��>�a�y�wS�D�Ww��׫����`��џ���^`C@(נ�>���!b�ٔP���`�F�IB%��F�ǳ9�sv4��A���n;n#�d6�ZrA�E���U�P1P�4*E,�����c��6l��u��!|�*�.}����^_��-:�/��dӇ������?���
�6�
�!��7�p�:=��f��W]��W̳DF;�b�__sF�X�d�����E��1��S���q2Z��Os�	�������gDq_}e\?貅޽��`���ju��'e$��Pe�Y	��X����ҋ�w�E^�5���M@�!�w��`܄(L�"���v�}���H=�l�Đ ,̸ivP�&��T�����;]Sz	�Н¾l��)	EE�!L�j��ЎK�X���lNv�����)B���8>[ɚ���Pl�l������i�6�w^SI�2�3s��lzR�*㤐�Pc���~��-֦5���"*0��g맏@�5!=� ���#�G��E*��^q%�cR��y��q��2+��5����@�L��7���[g�S|�"9����t���eV��f �IB��텎����I����
)!k\�
���Q��-��[�Uy��=;�䄜�x��cf ݁e�3A�1s݅w����}���F�5^�������$���	����d{U� �!�{`Lb���p��Z��e��EQ�dYh��#����\�Z�ˬ�ZJ��HT��0ur�{�9�&�TsZ> ��2lhE�r�#�ry��5�:��x<>��{���~���rz�1���%�|I2�C�
AT����	W#��M�ht�����[�$5���O8����_���	���7�w�e������@�ś]�K���p�^����:�( Ki���^N8�i������M���	�PA���~���kO�mkBi�47I{
���8���-�#ur�	
V���2�L
@��S�Bm�n�k�xs����P�[��=I���'����?�1PI�A^�/~�L�W�Sc?㕿����:�pv�ǭ+\
��U��˗�gt<+1 2�{�q��]�ĨS���Y������d��磸���9�Ч�7[^D��l����m�t��Fl
ė�a�)f�4�>IBW��%h�Yg��Zh�	��P��7KH�3뎰9|����k1��*=�k�A�k	q'�c�2�#N-�;}����1��8쀩RBI����}jVC�a���Ŧ�l�N�^�o��;�<*Vَ���dq�H�94y�k�mS����H���+�G/x^������[u�j�{yR��~�I<����3���J敬}�z���;R^���"���*��|ӌ�T�����4�\+T
u�I��$a�4�cJ��k�#'��V�a)�^��eևQ�9*����͛�$Z�)���b
��`W��5�w��!��i[��nM:���M*���ʒ��g��-��$�a*�1�6����a��g]&��$0I���<�rJ����B�{��u�3eZ3�]�j���ME%��z��t_τK���0�,D	��7"4��U4�P�}�V!<�����3�M۞�uWO��EbO����p��ʘ��i�N�6��ZX��P^j@��ת<jkgybQ8t[5��G�%�C�R��}��5Pv��\C��	�́i�MF�ZR &
N�J�1�^FV ��)�rt�����f�C���~�?�3xf����c�<:ZP�i�K����`/8݁{ӳ�7]4��nj���j�r���Ty�:�J5�ڈdb*�W���W�ܞޮϹ���fȧ��J-�8|���7�������S_%=ߛU��vߙ�P��o%0ZX��G�F���]_���݊�~@9X����\���ܦc.w�u�W����P���%�O��#9����Tq�}��32w�+V��]�qȖ��re��$,y*����a?�J�ŝe?��/�46J+ �):=�;�]h�b�Hpx�Q~�&��k.!N���=�%|����g'-@h	�l|�4� ~j�'��#9O�#�����{���H�b a�l�	Q(��/d>ѮՉ��,~f*�c�M3��馛E��ֿ�|O��	H��M�n��V��<W�p�>NW���	�	�z5���g�,�~���/�ʑm�Q�̶6��r :�jK�Ί�l:F.����\T��o��q����)CE���XZM8�0ڻYΖ������4�,�߼�|ݴ�;��ˎ�+1kjU/���?N�]�[�<m
5�8T�����ښ$�d�p@�z	1���
����BW՛����YI���=��?,6�d(u������C�S��31н߉�m�A��g�t��Jp?�Z8��1W�3��T�Tq>�V��بn�>+�߼I\�	��7�9��?�F�`M��A�i�@�10"��݇�Q�M��W��k�O�\z���མ<�O���8�_��W����EH|��%!�@�svg����_�΀��Q�V�BZ6]S��lN��1p)��W@ӏT���==�|�z�yW�����99�l�P�RC3��%,uK�)��_"8�v��e�.��9�x갼�ʁ᠁���a�9�4��z�T� ޻��B�
V�f��PH��= �O��t�J;[��h��e��5��
2" ��jRʁ��PkD�Q/�kƬ73�p)��9�=�E�j-�16���nr�-h�����H�C�9�*d��c)��~�R�t&�@���\G��J�FR6�!2�l:*�~���]�e����_�ѓ��뻐����M��a̚� �z��F�Г؊��a00]���ߨ2���q�IJ�.+�b[.:'2�Q���6U�s�LsQ�Ǚ����d�"���1�pR�����]�X�Xˆ�.�w7N86��]g��a=V���r4�!$��	�4��sW��_*ZLYf���|s���UyV5_���C�TMj��¿�5ak�ߟAGA��~��+r$l�~��m��ۑ�u�:_�MD.��@�C8�̚�M�e�}��q5����a_S�f�G4�R
l������}%���c��~�}<�nYvrD�H@|b��Un��2��$���H��@���Ey��9�%�:��Q'� ��넨y�L(�/V�%3��{����(��y�mGو�9@�H���<#<���/R'N?bO�����6(3`9#��'
�d	"h��9ܬ)�����"_�r�A9�Dk��GS�I��-�lb~���Ğf�?斡@�Ŝ��x]�l2o�-�"����;�Q��W���!���WWzY�C{P=��ia&�V+0g������NǄ*�P�j� �[��qR��z��i�x$�5�y<��q�LJ(t53�R0!)���̓�����"�Q�s	Hs ̆�ǣ�\�V2?�{��X,��R�ԁ5�����l�E� p��4�F/`pT%�����Xl�,��ӄɭ��S'�|�_U�#�����j�Hr�%;�MO�j�I$�vC�J4Jz��,mD,LC��ٹ�^*'��<	ū >����4��N/�^ti5l�M��>��+l��y-����YM ��'�%j�s_$�UlR!�;i�6y������$-t�wE����/�V�BJ�n��z� �JX>r���o��3O��X�-nkzPs��@���6j�� Yn�������&��cm��jdE!��7+5��^i=��N},ac�{���:O%�W�J�
�����bSȃW��8�#1�Km�?�4��k�G��>���}wv��_c�-[i���l#34�G������i=���eT��W��i@r��@{jv�`��Q#62X�_]~�]�XQ�@�2=�VFĕ��ޭ�M� �U�uWSf����l�b%-~ ޓA.����5��7��K�DYV��N�>V����p�`�!�$�Ѯ��:?����r��#'�2��CuL�� ��b�K}�|�#�lt^DcB�Ҽ6,-9��ftr9��ɓ�)/�U8&��j����gF1��;ݲZ���o��� ��0y%��%P��y�>��@�|0��~ϱ�6�e㯵mX$�V�!�ڹ���z���w�8T�.��绍���aPɠ�+�<�����&��82z��e���ٳt2�*�@sR������"�K���2�wK�?��V��@��}(;��X���Ip���tU['d��<7��z�be4�v���Z�Z� �o�R�׊�ݹ�[/���aI��1L�:-��`��W�@j��&��r��������q�K/���ҡd�z?�8�����i��yul2�/�����"f��e!h��9#�q�(�q�Ϥ#��=�	:Qܕ�/e0���G��=oNl��iK�k��H�r.#떸A���&DϪ:.�)>��6�n��Z�߮�Hv!S�n���e���A�;z�Ҟ������
��2m}�O�X�pFm���.d��:�4 ;�(�9}[�@Y�Ո�Z����n�b�-�f�����@p�+��b�v5�������9$yC�a�@����%.+ ��C�k�-��v��D������ N�F}��rŁA~���ė��7��2�|,~v46����؊�Ds�xΉ��+�I��"�Nz�2�����f ��i�2���̛B�<@�<�#�����ə6U�@;g�+;�,~mRΪx��&�u%IikŦ�8�	���o(�VgTd�C��'7$-3���e+MpL�XI󄁠�
K�]��_���yx2�\n�p��7�����	Pl�cc�c�P���=�ُ��D%w{'�i(f�L���.����YF=��ܮ؆}����G ��l&o��t��Q����:匿�z�0��Z�w�v5�P��R�	_�������{t�R��?�Á����#��n��������$�X�)5E'����f&y>Ӗ�a0f�����vKq�5ħE�B�	Ը�k���k_t��Ӳh}t��I�{�����e	�4�N��{�;-�\�1���s�9�1��8��@o>�y![9��H�Yǝ�ߗ�P���`�3Y�+V!����	�
Nx��4ƢqyM4$���ka 7kN��^wtq0���]�u�����I"A�a�����{��\U Ṑ��Ų�0{�F6�9�˰a�"	�&� $z|$�K@X�̂�ٶ=����/ruA,a�P�G 3Ͽ�c��y��M�H[�����'�������t�4�!j�b����@ĢKP̀��w5������\�,�[Ժ���&��Z�I�'T�K�iKN�ŝx��1��Dֻu��@[*x�I^	q�X�b���ywFb$�3)@W]R	V3�|��R��gPvTʦ�W�P�%�6H�1�|9��~^{�&;g�|����+�{�~��M��r�4k�|��{À�K��"]e!K�K/�m+ۺ���A�N��{��g,������d�&���:46��њHJ#�ua?��r����;�훾��];f���b�d�tl%#�=�yc��;�R'�=T(��u��Ș��r��b;0}BK=c2/4�u�f��:nB1�ܐ�:����ŚQ�B琅g�3\��pںu�f�k���:�,D�N����+�ƻ%B�Si9
tĽQ�#�W�O�P�������SUQoa�勋�R���D�r��+
|�9�s��e߸��T3ƹe �$���&�� �
)��z ��r�p�b�����#l�=�`ə5+#|��II#�B<>��i�|�T�����1����`���y��b�i� ctxfF�Uc��ǧB��P2$�._�9�_z'B�H2\�̞+�9�G����Y[B2�Zӊ<�8TV�u��+Pӏ6@��������{E:�:xg�#C�HPp������1؂�72�����r	k.	���n����C5x��n�y�K���]���H#�,�Q���
nw�����hj?�0:[uͫa�i��u�������;v$Z	ᄠҺ�g���L�}��݈e�hF��ݫr	ΓJ�z���=�`�����;&E��1S s���2_�(����8�MX������O�&�DĻ be�O&�M�sV�PI��X��K&l=ާa���V�;��(L�*{HQ
�8��jn�z���F�( �\����u8�ۭ�X����{BӡR���������Ŗ�fN_n �vl�J�����Pt�B�k9b���t��*�wCR�eGC�/!$\��Ȍy���7_t��s��ӌ�L?�L%𬦵
nĎ���.^xl��� 	�S����fΕ�l,���-E���=4���}J?���\46VI��ah�㩕C[��qa���{D�vFmā���<5��+��v��ݏ}�Z��~j�b�p%42��r���/iwJ5���/\���RjO��K�6>�"�,X�is�G2O���끐2��\���0@�\B���uh�4d)�f�)�i��kk�J��E�B�MvR�x���R��q�@�Nz�/���v�z�kEC�;m(��sv�Lxs�����*֎��ʗ�g�//�*�$��o���ny���?n���h�c�Eڣ��YiC��xPW��b��^u~���7�������G�q>4B���@�\^��
��7��e��c��P��ܯo�g�F��^�G�/�q�H
��[~���/�ᣤ�~�[&!�%��bt���G���h���星�T�C��=����+W��4�v����s����۳h�_Ѝ"�1��(G���u����b������0���	��l1"�2��v������&���Dr�3�ِ��PF'�����uufP�I���]��D�>�6��n�Sa>W��퇲W�M��ޕ�����^�"F�>�%F���iyt�
��3�e��`<�%�J`AsS�S1+� ���}�9�d�d�)VŜS�^Z}C������v�S:􄪚�~js��X��QΛ�g��2�Ʌ�� ��󴽫^c������M@�u�9?4ǻ�6T��"N�}��*+S@��Ɖ����nN1}BU�V��me<kK��v���-C���w���K��Z~�'O�\��p#}�uD�q�\ԟ|�oLnE%c���ѕ�:FriČ|�����$�6��9�"!�p��Q �Uvx��}�O�y��9DQ�ߚ��Q;�W�EҢ�&:_ܚ��]���~г���b�&�H�*J��;z�#F�'!�4�S�OLx��&ٲ��
��fZ�E��E�y�c��&s��#J���/C�郼I�6�+�2�i6�蛄J�ڑ�,{��~z҄O��H��P2&%�u��Y�<]ù���x\=�dk�(,�!(dfAR��Bl�mr���) OH��vg�M��u�{�K�lԈr({
v�m�x���L#'߁�'��pO\���"F�$��z��.Z$��>\����@�ɩ�͇���������-�OJ���Y3~k���KY��DЯ���*WE�\c~��W�b���C#�sP��[�_�	9" nݵ#��AeUh���5�yT1~5���o� AȄ1���t�n�v�;��?��ݷ�>E�iv��kBё|�~��rM=��[l��� )�[��[����'%e%�z�!2:��t��t��U[�h{���&��Ll}Ka���Z�m��@A��X�0�l U�8�Q0��.�F\�%�{"��޺2��F@�p�U�����&�`��=�^�x�pu%���ot-B���IK�����B@ќ�S#���I�_�D��5��Z'�p-�M	��څ��'���������\0m2;������L�|����tpg�x^��GPEa�R+��_��ćX*�~��5��� �#�we'_fp�[�4����Ub����M�=��R�nv�H��2��9Kf�>p���fd'�o"�0U~8_��O6I~���ߊo���`���� ��n �^�|��{vvDJ{,���}P{6�:�N����
�\�p�Y˝Z5��V[�?�D��3�نV��lW�D�l�׸}@;�}����}��%##�H<q�Z���m��U���G��M)Ii4����V!�s-��ܚ�����A%��.(ioο�����K�)]�Mv��U*�W�"_Ba�~��Ⱥ�K�L��	�}�Z�����_�#�S�6i��$p�Y�<4��4x��.y&���Ǳk)���p&,�"լ��)��mx�ɗl����q7����`!�ߩ`�F�SV����lօKgM\�?a9��"?�3�!�H�Jݠ:A��]J�ǎh�K�v��.e"��B�Zikխ��D$�v�^BT^�7J9Q�Ϥ�cq���/U9�g�����n&��e��5�������9��V�R��,��Tx?3"�D�{�o��#%3�4���
*^�(2�&{	���������חE��h)�m	�Xe��_G]�±��Lq�A�R���tӪ����Be�������D&ֹY)^r]Ɓ�ui.�9m��凓\�E��qN2��T�Q�!�VWu/'���ڿd��۶���KPw"*�����y1��%�&%��,OE݂:�kK�t�چTH��6ڇDӪ�o�"{��η���(����)��W�N�9v�ۍ����o����|������FR ���{�a���r{F=_���V�F�u�\Y����=ヱ��}���O�&{�j�zN�����WI���7S7�����9^��ݲLx���N������=*�Cc���r[��'R����Ӗ�Q�8�s��_$�2�<$��<N���f<j5'����cn�%�H����T��U�S~y���0r�|�${���(�gW��|FA��o��N/)���|J�k*a�x����ٷb��۬�4HSS	�X�Y�18��ݍQ��Z�@V�Khi�&aO���3U|���t��J�v��Ƌ@B��݀�goq��?�#Sj��I`�*���c�����T��I�C~"�t�z�����X"���n\�ߨ��^��r�u��lӭly�aȵ"�)X(���H�G���lA}���IQ9v�?�gY叮������Jb�4��E�'�92e6>m����ǹ�0�U<b��'����	�^��~�HV3�GB|!9���V�ȧ�A��5�~Gra!X��m���K���a�_�+Uv����̓R-o��H�9�?�z�K�T�ĝa겒��\���U��a����yf=���u5����0P�Ų֡�;U�kNq;��jv��� �.WL���^�9�Aq� ]0���Ԏ��$ۅ!���%�i��������A�����y�!}� �y�l^pf��%	g�e�%���ؖ�=��b�R�S�V��tOD�K�j4r톂:�\��3�Y�u��w�8ylL,�����V�8]�ƣ}Z��U�D$�	U�UC��h9a���Pͺ6��ch[=�G	�;�� S��`$@�����s,u婒K�̉|`��3��}�!Îq��_���F%�~�{@���{�f�Y�|u���t����J6��*�H��	Qٗx�]�����8$���~h<�-���x�R��I5���lP�B�z�=-߼F���5R!f��ài���8=��ԆE��3��3����t�3��\ ��w��z��cIjv7��$FBJ N�>�j��gM��ԸFSR�U�	�Qm��X�û�iκ��x�I����L�:�'�E��E�g]�<��W�ʦ����xON�E͠�@ 짎>_�|�2�Vkp��ƒ��Te�{�dy���̯���b�N�����>Ӌ`\�Ap/�֖�s^A��e>w�Ca	?rBY�#&����5B3��r���1����MzN'��U�����\ښ�J�wlUH̿�ד�'3��V��.�J����:��S�K����mυ�JlÑ\���	e��	���AP�|&�$�;0^�8P����l묶)�+
D �m-�= ���"��G%x�MR��G�x kN��"-m�5�Όl$�Ժ���e�������/���
=NfB�.���e8�mmlm��Jc���pz8 x6������j4�(Zgs���DL�ժ�#1[�t�3�Ɣ����!4Z�|��l%2����x�u�K^*�ɠ�#����e�c`��z�������_sQ�ISXf��*����A�K�iI+�m�4kc�y��t�М�IW����$���c;����<���?��GҤ?S`�w9�V4!����8ݝ��P�T;kH���,ͱ�R
�|�`//e��傐h��!�䜽[�]z�w�z�DI��2������YL�f��bp�J�9������p����f�F��(҅0r]78e���V���E�Uܾ��F��|`��I�vwW������qmn`�Q�B4� �8�Th���������TM��Օ�ѠT��w��4�6B4Y�>���k|%qO�	=�{`��Y�P
��Û,2�Fv�m ^U��Ea�b�^c�柳�z�%E>��ө��9f�}���;�U�!��>���$�_Е�i����bG�����̍��Vn��p`�H/�'��Z܅��\e@?~5�X���jX:���[&;���]1��>ر�2�J��(�T��m�\Q<M4J�8m�oZ[L'��3Zi���8�� "�m�Մ�Eh)��^�<7�Us�S�"�����D{y���ɳ6
��)����.�s;���?���P��ߞ��b:o�[�)H�5�~���Ԍ��(����%n��{nŋ��)Y<�^���`���/s���n��1Zh8C.u�m݄V�ʥ�U�H������ߺu~�p�@�|�9�ϛ�	!���&�u�:h[���R�L~a��ri��r�.�ls��2$��l������G�:�k��_
�)��q	� �PPR)i�;���?�x( ��Y0���3��&p�Y���B����\�݅���@�YraV�5!�f���s�}�a��p�������OpI�@ ����$¾u�����X�⹝�#�wC�C���U��z#nO��i8���QL;Z�c��0ds��ea(�s�.��;3��i�SP� �d�T.;��4�s�}�w��@^�F2İp/�_d���O�u3���?E<5οo��W#'�̱I�U�Q"�t�J��ؠ�1�ddg��U� ��~hA�p�`���.�K,��l�J��[��@GoG �"�Yt׆���&����,5O#N�;D!n�p��i^�,B����<u�����r����T9���'X?TmQ�!�dJ�̀U"1��š��L��G4�pHn��A4�*�8���E�@���k�Ŭ���l�tj �7 #O�Z7��#���_ ��[��*J��j�	C4J��	�A����h���^$���M�߶v����\ �l�S��)��̈������t��T��2+�D�ڿ��{��\g&�Si����g2�E�{j��6j����C�m�x�OGpCz��R�PdLbNu�\�Ӎ�������Fh���B�^��T1�*�i˫�/A}c{�t]b�Y�l�8kرx�?a�^��sÔ�1��9�a�$]����"~����~$��{��i��G5��z�ƥ_|�,:���A�0F_���F�8.Z+sXfB������yZ���Lp��	��o}��:<I0�WS��cc���'�����
�^8�oȁ�[��II�P���汅�a�rTS���-Oٖk!�kЎ(�����S���������n������Y[��^C�h�n���>��]�0�}��4�s9W.BO�u�����c�sG1�{���w����9\���j'�o��\�V�Yn�C��Z������R������0ڶ���+�UR��	,w�d�(�l����%Z�(o��vj�!�24���_��ggG�����+�;�:�)sa��Ȗ��,��Ԁ�oM���ܼ�E��?8�y���s6���HɦB.K���y�a�i�5�wܜ��گ�v�	)�5���v��܀A�����6����(���O�@�ф�7���Z<�S�����m��.mwVL�ǈ��	�:�p#ԆD��<q'��`3�K͡��/��x�3��^��u־!y{L�5�
`;��'Y������3�7����	���;0Fh�g��e�'�#�k������Z��`����O���lF9z��L(����$�.�0
��7��+�S�k^?҅�Ų�X��%��'����)p9ԝ�o+]�<g΢`���j�8xny�ZDڸҞïy��д$�C޽8�bIQ�!T_!�@���ZH������'M�Y�tB{�=l�@��|a�����,�4��q�[��{�z�������E�0����U���sXU�����sP���G"䒃!���(ˏPlh%�����2�/��0��_P�5��L���B�g�~�� �D�G�:ܫ���%�(e�b��+��� �u	���/������!>�&����n�nvĜTK�D݁y{�����MR9�}nՠ��]���+?ΖؗQ�Ӕ�e~���RS�*�gu��y�����I{�ÛA��c�<�U���c�i3�Lof����� W��K]Z��`2�V���,����{��,�L
���p��c�u8�]���V����i�+��:gP���LYX��zҿ`|����a�W#oM=���S�a����mBK'�r����[w�`�,�������������m�2�o\1"=�!��L�c�>`]�QT-p5(�n�;GL�Pt��*�r��[pZ�;�Mu��o�f�\1�XW���S?�Z���W�c�J�J�m��@�A�近��U��
nf�C��kep���,�-3�F?��i���Hm�0��^r�⯚o`��2?�O����YNĎ�tsC$��fIg��yR`m�6�D�U���J�*�*Q�̂��)S��F�"<���p�Xkj��?���ꋉ*S$et^�� ]�H������|�O8��/��m�/���0#�ٛ-A��鈸}���F��g��S?$Jٔ���G����+,����RB}�Ĩ�����S�@ޯGidXݕ�D�'� �� 2o��y���~d�P!��P��z�N��z���b�����l�ܸ�_�Mu����	�c�.��C(�������N�*jl�[�exQ>�:���fB��/6M���t�M�=����\�m�E��X�j���n��U�`�N�eG
�k�)Wo)�Bs���h!���x�:Ϋ����G��R8O�]||Q��vq��C����0���P��%!v ��*J��&�PV٧|��(����0U����-������E��2Y�~,+���6NA��p+_߫����<t�#Z5��?���C9�]ޑ��I��C��k�����7��b�TK����P�FDD��4��)�$�����*���G>�ל�=J����%RI#��=

i��C�8��!��XD���5�ϝ4H��w��r��"⠋v��nە{��}謦�g�-&����؁z�Em|>i�u��sa�R 	K6cG���O��b)2���]�l�3�ȭF�o��0_���G7��#X�@$�9��Y
�+�U�F�?[��	&����G��n���<�ڵ�q�yZ�V���Մw~�l�&�6�r���mxΏ�M����$a�Ξ_ŸK����_�S"����t&7�4'�1y#Yl�T�T�s����N��Z��sI(~>os�a���:�q��-�^j��9��j���<������M�������d#�Nح�W�0�U�Rgnx���?�N�+>�_ ZΐE$�׺j��	gbf$xR0�K9	��2JG�l��q����P���O�lD�83\�7��l�'t�Sك2��;�F�T�|G!���$I��F�������6����V|&�[�E���R�&�͟�b�A2���c=Ř��4L��z�F�!�5�F1�43��Ɏ��fm��D�N7��`š ~Zu�k�4
�3q�6��;.|
k}�N�{�����pMN�,�iVn�.������\-���!�z�Q�U@�f���m�P��cH-��f5Ip�y���ܦ��
�5�-CvҼ��w`AU�*?k���c���k]z?���RZ�iy�_N=�ʵ�3�SHQ� �v��	�*ƃ,��戭;���c��]�*����-v�n���#�/�V����-�d}�ɋD/�-&K��A�;*��43��b����M�BCݲ�����hO9�)3^|����:�~/�j�O�,��A�I�Jf���r���2��a��P�,��c�x4ߤ�ܰ���ӻ��s�/�~kwR@[wz̜���ٝ�ؔ+�c$L ��COJgd)�(����=;QLn��װ]�WSn�s>���u�]�p���"Y8T�6��B�J��w�˻�����l^/����1��i�w���b�XO�rf��0<罺W����qt"�l3�
»:}�ۜ@
^�c�<�SRW�|�I����ɮ��6=	����XZ |c$�)h�S�xJ~�c&��!E{��j���})%{�rn��;,0�T���Z(�,)h	��s��!����=�&0t����C`c���xQG#41���|�M�����4�R@�S)w��أ���*�P��y�Ѻn$��C�^��w�`$�Z�1�5w�,�$�XoA 6��;����[��_9��"ʾ#	miτEc�4b�_�(Q���h�mX	���%!�w�)�K��֓�?�g��6�q�YP��P��#���L�(/_��,�U�����,Y�Ύ��5�зf���g���J�(x�������P��j\�ڽN�<vF�}�FTs\��y�\�����{Z���綣C4�L���>�(ڷU��l���b���\���UR.�AT��������n43�6�7��"a���s����Z�Y�����fF������w���!�[����-���r���,!�
�5!��{��(^�
C���;Gq�V?�[���K�0��S��oF��Q����p9�{�=Hx�? �:�aq�6Q""���u���0!F�[�*e�Qn$�qQ�X�/B��a뗗2�.f��9O�-,��VT�~`u�KK�@.��(��]��;c"Ved�����s�.��D��ʕ�={j/�n��ˌ/3aA���Y,Җ�ŭ<���Ew��ж��)�l�/���)���E�	���}B��Q�f9�Ȱ�"@�z#�SJ��n��(zӸ���P=gs���(=���Ό5@�t�]���P�3���l�E�F��٘*���N�����ʗ�۶A�N���"}�Nw	�]�ϥH�'�I���&�\�A7ż��i�� �m�aޘj�Z8j��&��'4�q$[�"��& V�G;W�Ğ�5��_8fG�>;>���hmr�*�p��Ig��sw�9�k���6��A�8�����]!Xnq$���ݰm��^a����r�+�e{�d���Jҗ�a*��;,�B�l�;� �JD�C�J�����W�`��''X����¦೾�̓�	�N<����퀽��{�\��⚺���.f�d���zq\�#��z�)�%[��¨���4��s��� �]�u^�ڗوpP3)K'>`d��f<-�T K��Z�!H�����N�����l
/���"0�R��F��.}5e�s�X�Y=��c܊8�v�G�������-�[١щimP��AI���5T�j��1�71"�l_���ԙ����� �2��7n���|	~X��H[g=$?�"�Y��������#�&��$��ϗ�X�}�/d��ȷ�>:� ��wg��"���\1�~{��(�'<�Y�L!�id<ŉ�Xsf����HC��!���{}j��m�j��2VۢP�I� C"Ļ�Tw8-^��^T�=�O�0��u��u��'����Z�J:[�Nۥ9_�ZAA�.Ri�D���'�6�Ta]�/OH�L���d���$�BeY<V�]��b\H��#$t}*L���Sć���u��"V!��Y|'�,��U�o�C���
�lU��r'�q�i��0��:Ɯb�)�U��Жy���G���Q�m���$	����tr5��)g)��t^9M3^�p��U	W.^��{p�*�%�x�{笜�^}U���� G��2��%��H��-'���C)�J�c�.��Y�o>��Tbad�S����%'��`���e��l8wmI���]��5�h�P����3.����+tU>ʴ��2'�@tӇț���|�#��U�J �/�6�5����?���l��c��/NH@�a)K���ʠј/+<J�g?e0�bE0u�B�7���ڱ�/�5Rde^���<1��l�:آO��E�(��+_�Q��� �U���=%h\�Tބ�v���ߣU�d������(.�m���	�A�f��Q��w�eHq4�ev1,S;�u�U�� �
ݯ�2��DjS�W�KE3�����<��l�U�7�<��\���(	mB#�Rw�E�Fi��,�Fi�ߔB�F�\�AP�&; ��構�^�K��gkX9�s�1K��̍5c�8��9`/9��*'�.��	�(��R:���(I��){�|V҉��B�i�a�@$qrĶC3 ā��8�u]�x>���k$���$
�k��]�4t9�e�P$&	A�����7�*V��T�H�X��2놱���#��e!*���>~��Zui�J'Q�JY9^g�焻��>�E�`�������xD,��7C\QDI��9ְ����"r�i�}���]݄7�uJ��{�vճ������&^��~��ΞP�i<f�Z�&5���5:�~j��|A�8f�Cv�eEj�O���cMsG��#*L�k�N��p���'�re'p8ސ$]]}��];�t����'�-�C�r��w��Ђ`����5����7D��[��Cq�<�Sj�05��ēj�x4�i���>Aͮ�\�@��|�"��Q��.Vn��q8@51�jh4,+��Xe����<H��R�Ҥ&p���u�Q�	�μ�`��8V��d��bF7D�J��]�+�_r����БU������Z����B��W��=:N�zQcJZ��'�v)�CpvlH2�K�¨��p�I����䢖|܉2�j*vۇ��&�9�����N�C���Έv�C���L��S����ζ\ؙ�)�M�B"8�!�H�km��T�����]6�RR��D�R��P�`����?���� k`=�(�����1"?�k	�AXlcnn}�.��l�X�1��ؐ��!J�H&y��ދ�bt�@>��/��\��lj����M�n�l��H�Li��
8sV+�4�6FQ鎜�.+@�����`�_k@b���4��|�3lS�F����ȿV����93��we2zG��v=�-�?�6AA
a�R��}�1��6�Zή�Ы���Zca�Pv�|< ��#�_CBB����KIX���=GrV�D���-$B����V8o�7UJ*T��j\�3�r�N�]�A,��ّ������I
�`���"l�ٰ��Z��O,v�4?�U�.��I�[��U�1���������e1�ìߪ`$������&:,x�КŎԑ��R;����ᄆ�������s3O��\��u�;����v^�U"%/ΐγ��P�T�g��Pj5j��M�#lU�J�Rs�hQɯp�0��\(8ַ_���^f��ݽr|��hD�r�烴��Ĵ�w��/�,����>�磔��Ase�E�"�������ű6�`r���v#.�Y�R�CC�ͥ�r��%l��s)K(�:��C�����uΫ�ư�6��7���}��Q���Z��ρ���@��zXN����_���_Y['d?���,s�ʉ��w(P*��Ḳ�L�}Z}U}��B�5B��P+go���1>�����N)M��2ͧ�^����V_צ��\���'K�۽���[��A����-�%=l�.�S�dPr���#(g�G�NK��t+�YS��%���d,�G�:�؎� �J1n�8�e��ǺZtri���Pӆ��?B���~���S��Hㅘn�4�<��0��(�;ؼ�H�i���a@Fа�D���Q���n�?o��7%+}�������y�x�F�(����T�n���P$��
��X'�ip�[2����&���}�:T�R�ʁ���?/C6�mhEpB�縀� =��?Sy�N�,���T�a�T@�`�!��3���l��:��D��t~��?�U˿	RO������G�����$�(n�[�r�� ��y/ϒ�������^��8��.Y�g��z�!���.۹� Juɥ�zq(��0��!�����l�����υ�7+N�`�T�6���"��Ss��G}�oH�^�ض��l1���S�@��^d��Q��[��দ�=�J�
hT���	��azH������l�n��;���h���`.��i{�K�'�#�n~�`��@]�'bx�5�,C ����NՏC�-sؖx�?h+%9�̂��������y8��#���!������,��X�>O��bŕF����dϒy��
�a 	�i����^����ٚL��H�V/x��t^�QJ��J�>P��G
�ʲ:C�0.+9рQ"/z#+�L�	����%�is>�����6	���q"ՔhY?�%�3&2��\j�� R�ҦГ&\�J�5q��f��	i֪.�Gd���%C����d'R_r� ��G/��(%Ȱ�!,�I�ש@�:�x��T��ɽeSЍ��ڊ��+ʴ�-I�ɍ��|!��:P��3�|Ҕ�tִ���{���<����a,�� ����76�H��Ō�挴�pD�&8W΅ؘm��I�(�,Q�����3�e���MA�L��0ٱY�Q	�>����y����=�
ݘ_}񅇨��*��9�S��Akc~���e���!%���73�@��QY(���D}�YbF��(C�I��)�!K_vցk�,I��b�Q�~3]B�6��rʞ{���W1Љ��`�`����_}�DB��.���ņ�8!;�S��k9@�~>-殕��FqW�N�3�����Z ��La�]<����kJ��m��J�O���R����fXw�j�du,tt����X����=.Ҳ�����H�C��[�|+%����-�:��bX�,���|}������M��qP�P��ߢbZ�!MK��7`��g�0T����j�(����Z!C���}�=z�O%�RV�d���}&�� �k�"�>���k*8U��88�����7K�2G��[>�y���^,U:�x�)��$�D��m4��m��]Ӯ�yi<*׌)=V�#mm'Gی�5iyll%Uw�K���B�����Ot���c�O�"��S{�k��pK��ڴl'*��Ae�*�V��2$K,+/H�/��罶1؁��N�	�$�Bxj2�#k2]�8!DX�p�-B��Gp6 a�m�KzH���#|̖��1;_����M�bE���9�!��a<o�&:щ��Z8������ �Z�Y0m/P�uTK~
G':+/�^��V��T=${(p0�[M�#�J�rk���嬁R&�K�賞����f}�ql�Gl���[z�j�> ��.P�-u�������%�~^��{T�X<Hs����%b\�t��n	���^�%�����]�8��<pf��
���)Ð.+����*Ni��0�Mo1�����T�|��.��h��D=X��& >ϥ
f�'����ҘﱔN�����޶S��Y�m$��C�&��:@4���{So�q��ք�����̯�����m� ��wƃ�4�m���ҭ�H"� +s�T����ܷ������Ӹ�,����*ۘH����!��r�_�2������R]�_ ����\�!�༫O�t񚬗��=���m19C��_�^x��)z�j����%��oѡ`�.�,+ '�	��޻ή�9��b�#��J���[c�N(�=$��V"x��먘:����qK�1�q�o?��V�]ӫ����?�S8I�/��0}j�l����Жِ0�%�cN�4���oA��X��fM֊�f1`Qz$�3] )�,	���a�Щ<#4����@�؅�v�u�Ӽ�����>�VRrl�I�kx-�ʹl�Є,�H�r���4�1���.S���h&���=zm��;��>Ѣ�UB�����+�Hi����F��!���2	9ѐs�v���ł���l9�L�����_�K֟�ϣ�2�9)�K� �QB�pS-v
No�L�K�)��*��̦SG4f�
�  �z`C)"����6˞���[��x#�VV^:}�y�oVcXȾ�����M�i׋�N`��<����튬ع|�%�B:#P�6)Uc5{ltx9�
_Xƌ�φ)�P��ɻk���b�k!��O�m���d���26��딲=fT>Z�"H FP(�}8����!0�!c�{D�L0��L:�k6�d
zT���-����3����,k��Z�n�a�����j��"��s(��!�0m(�_�mCؚ�k��[�dh�����ڿ�����=�}g�:ZoqHzl~Y�g�h�&�qA�3�t��"J��ibF���s�GQ�~�1�n��D���k�o�P S[͸0�M-FS5V�כ��cy�Q�%!7�FS������JJ��ь{0�z��'���AwG[)l�]⥰�����P^�np��39��.������	N�n�B�$��ܞ���}S89�γd����t^�e)N��淯v'�uk�&�r�K6��Q�kz4\ɽ��<civ��k.h�IE3��G�n�i�x�տՋh���{+�wڨ�31�b��u�zq�-�<|L$�E1���×ե�i�ڱ���CE^��i�z7��%rО��������k"��3���j~gQ�4�S�w~�~�Zc2�ϟk��꺝e�M�*�a	)S�r9�G� 6��q�N���X��l��p,��)V�o�����q��� 7���
U���s���f\����ti	�2��x����U�Tcea��GA�PzS2��k�h��lp��ď��*�69�/Rج[���,le���?��7x�J� �NAp�;�c��"��p�A�z���򿁌���Uix��>f)�?��D�܌ۅ�� �
s�@`���n�b��|/�����q�pl�o�Q����P`���Dg,��"�ߍH�b���3"��7�d��RL�a�����rn���zq���1G����O�@�S��ਫ��Ih]dFa��mZ=�=k�խ��â�Q�W04)=}�n'�~�3'�å���;��-"�M\Wv�=�(�9��a�l��)G8п�%�u�2Pö:5@G�F��E�W�qVbӮo�g���ݰQ���~��nR�*��	R ���A57I��3l���>�g�
���QP!?s�̫ట�x�x��?���<���u׸5�2X_�U,~N.�q�l�fQ��F�n�9w{�Gb��@��
If4�#łK��6UO�3k�m�1沈�_>\؇��5���>�B$����ӯל?��jU��^�)�T����pș���.` ~�"���k�ڲV��PF��5IҀ��%��UuF28#�xrqa��H'nv=���/h��a�N�I���&��"�<V�]�I�x:E�;�Ƶ\�FY+~���gh�!d��̵��T��D�{�wn�%h�l�쀉L����!�Ɯ����`������3�R<�QQΩC���{�j+V��=rq��X�ECf&+�ׄ�)[��Td�风2-�����݁���L8�-V�&��#l���JC�R#������'-��ߤ��8�����MD��˴��ȷ��Z��Wlq�G`����� �)�i��YFL�	.�U���~h��Ad�o/A�-�0S!%ЧVw �	~����O$�-���`W�*Q	킪���O�����g��{��*�B�#{s��$���:X:_���>p�m��4+��$��Bp��ە�M�G+����Zta0�+	�WJTR�ȝ�C��V@-�%+���w� x#�A<��O�P����>=n������T<H�Љ�T�nbx�W���HXx��U�9_Tz��Ft\*����J�
�I��a4�Ce+48�+-���#����_@D��^�H�ׇ!����R�:���)b�ia�6����)\���<DC�^���>��\C���<#�ӌ������Q0��ڋ��0�I��:2�GR����%+�O�,�9����P��;��6Z�(�I���e`��>����U�J�o���
Y�߇O뗳ST�y�R4	>m���r�r�d"L\��U)f�	���!Y����2$����9(����Z2�?�M�)2�Q�<ٳ݁eVF��/Ԭ�V�b�Q+w�����-TR�t?D�3*����"�"�FpZ;'Ǝ����Z7�i� c�s�H�W����J���j�S�&����@[dV]�;��V�:!D��wUnƜ����[������<xcӱ�#c
ܻ�
����G3! �e��ω��f�<��;Q�H,�ǲR������Pk�p�F����q�8G:A���$Ǎ��3�K(E�u�~��jV^�$��zH1 A!E��,���}�|���bv�����'�*�"w��<P���_�Q�>[�o�Ӻ!����ڴE�8�O�tg�����gl,�� oK���r�����w�or�d�E���Mi�E��#�"��u��Q��4i:�KFa{��qH��}���-��]>��Ȫ��s��/�,�eH2������ ����
�	�M+Ʀl2+� ��/��L�Ǩg����]W���-�&b5�p8�@Db6��]t��p�/8�`7O�D��0ߛ�w
������]��p���mʣ$X��,�i�|ҫ�?�3B�0
�X�-��!s��V���_���b�	AIӥ=�M}#^u�(�wǘcSc	�(�bkf�s��&����?��s0܋�����)�|��uV�?���nն~�S�(�P!4xߧs?@ D֠��^�l�ϩ��7��g�n]
ט�[�{�`]����H��x�&�3�9��5��ūI�!ȫw�O���
7݂ͥ7�68��
m����z��~)]�d�� �R'ޘ��G�M`��&�]�C�J��=��E�Y&6)����+Ќ����q��5ּ�;�Ү	W��!7|(GyQ�A�gT�B������}"N��
	C=�RETXA��Q%�
�b�@tW����3���Ĵ��H�SQ�`�Y�^�15�V��d>O�H�ED#���|�6 F��\Ls�f�h�w�hP�Z�{z�ރ���j�"Rs�E��V�h$fyٲ˜k�2Q��]�C�mQ�D��@����[�t�ڼ��]��{�9�h���P`��S�TnA�h�)Gj����P�2�ET^>!s�@RJ���S9��9|�t>tE����y*KT
��Pr��'H��V	h�}��y0�[w����m�
��v�VM���ͨe)`q�q�A�Q}T'��_%װ�;a�~C^PI�2O��Q�ϳ9��_����s�|hq�]K5U�9��$Q����<}LJ@��U�n޶�\=;^ ���H`�|�"�G�Ւ:�v/��g{�z�v+��A�:n dҤS
��EyX�X��=y����z˘4z�Z�{�g���T��Fy�ǆ��JGE���5�V���w
o�A.m��/��$ѥ��V#_m���zG���qv��+ۦ���x�1�0%H��~q����7�ić[�sJ=�ې����:NU������c������<&@�a���y�Z�U���o}�������?09*�m�y����e��\��
�d�ғ�J2�F��f�\cN(���1= ��΍��C�}���d�o�� L{J�ڴo�IA����1��0��'z[]<q|�j���`~�ǔ�4Ye��գa���CZ7����5	�h�lk�d�*����p��?={	S�i_�6�/%b�J�-��*óS�����uKD��c{6��T��ё��8��?rӟ�]C��n|��5��$�m7�o/�f�in��,���ZL����A�����ܛV�Yu�{v^_�;�X���H��dz�ֲ�E:��dW���E֤��b�lb��+M��Y>E�n���D��Ͼ�d�?���pvg.�u������tl���ؕ�]�TyG����򈬱�Y�q4���I�"�L�hy+�� ��EY��:��Z�~���P� II���XA��B��x^A ��.q-��+l��ws�L9
����vc�n�+S�1���h\#&=���G:;U�φ:/gYn����f��F�]��(OTW�5�!Y�;�.(V��;�s���u���Ih�[?���
�#ĥ�wwQ=t�'��T����<���zMtP�GBU:���vE��h�4x�Qq����u�T��y�{5=����;|��\K,� q0X4��M	�׿��G�1�-�)�jet�c��$�c���ՑC7�Jk���$���@ظ��Rʫv>�����F*T���̑��H&��_ۈ�{_+���X�j�8�{S Oy7i!�*԰���m*Xn ?����P��������}��,ȊU��C�z!B���!�>��òh��Xg�3�'�O����W_�܊��*��c��	�v
�����y2�	!(�eJ���/IA֙+8]{5).�T�9t���bb�8� F��`�����Ns �Yh,��vx��a�%j���p�S�6��P.����Vo�+tq7!٭���E��
�A
q�T��͎w�9�I�^"2��Y#�?d��QF
t\��+���뫥l�����h�h�����A
�5�+}���ͱ;8��<-/�:5?��4���W`K��|:7,�їÃ��y�P��� RՂ?7y����ܨ/�,+��.EdVT�j�@�D ���o����G"�����86�&z�R\��ڮ�J�<Ge�b�/��}k{��n+��h9�0=��=�:������ַiɘ��4Q��b�W�RE;��UB˫����U|�h���B�˵��v޺�� ��HX;�P��j��?��*����$uP�����ph)ޓ`�I$�'H�z+�	�(
%}����PfՄ�ZT#�p-���FY��.�&��7��$�����n4�|_�L�l��*K��]��D$�.Y��w� 9�]KG�'��5�̥(������O���N�_��9�jή���أC@Wm?�f=t'/V�1��C6lvOq��䑑BX��)Jr"��ޜŻ����Y�f/Ey�	D3�?���F�sD��̻�#iE�ن$�DA!̛��S�!#��f�E�)zR�ۤ,��=�[
z�
�#������B����L[9����W�Bl��e�O�;���M��@U<�
�&�Hs[��{�V:�v�e{-Խ��|���Ҥ�Js��a��L\���.��1i4ؓx��6�$��5r����+��<�̙���Ux���d�b�gG�}<W��턁"�g.��ØQ��gB�ЀS���1BK^�}��^*�I��4'�.(���*@a�Sf�=�ۑ�{H&.�3`�VQ��&V(c�RI7�V��E�H�?�}�Paبn�V?�hy��u=����!�;$�t���z�qѥ+g��?#{\$��xVT�hN��]e�����+��1�����7���P� i9���69�
P�J���e���s��{(�z��K��ံ#�8�Q<�������yv���J�l�m��.r@Uhrx��>8!�Z\{�1��'�
[l���g�uՋ| L��G�A�x��z,r�t�;i@]D�as�}��{����Q��������c�)�'�4b�v���߲P�[<9�9�vS��I�y�x�2e�)t9|p�B�p��wmU�!^zc�2�p����8��4X��78�S���[5��(��m��$�p����@3u���o���	.�M��e	������1^��rn2�B1Jp��Ou��d�q��S߬�Nyc(!� �ŵ��^���Y�
6Y����HH���:�����}=?a%�R�'��V7�Y]��cr���ٸ�T9,�D	ϭ]Ɨ��*:�H%l��*?_���3��5�~��ۤ���� 2��ҝ&��D��V���4�9& ������6���9�뭧��c�&� �Xn4LؘE9�a�݉�;��Lw:3F+y��E�j0.1O�k]�'�ǒ�����n%?������.�tE&o��w������i�t+�	/:@fG�	>W��lb, m�1�G�V�T���y|+_�O���ƣN�H���X���u9ʍ�g󊈘
я�o��M}xs�h�V�Ó��q̳tJ}�6�F]7�Ri?�'5��S$=&��҇vʴ���#H,�
�7��ϛ4ȹ�ۂ�*<�Gc��n\*M�E��=�
{�H��Ӧu�T�®}�L5\EW!���8�\��y��,zȐ�e�5K:�+mס���=cB'�K��Z�d&I�p��`��\^	��������L��6<-?z�'�=1v6�7+��p]A�"�w無���o����:�H�.��9�]z�+�F4��Z@�=�T�a�
��[��
j��u���}6A�}%	�h�OCV��of�}X'1�s���W���cy�K~�^N���<�:�G8v�H���;� ��v���Y�2Tr�ؒ��ŝ'�03�3���M���U���`n�-�y��ͩO�3���#���� 7� ��o.[y+9��J���|�Ȟ�	($�����=� �Kpe�։I`x�=�"Z�����̓Y=�b���1��,'h`�%=`��˖T�_��k�,����Rz�Jۜv�X��kI�; �&���Zͯ#�������m�E ����0K�Es]�x*˂� $z��q�W��?����."������hI��v<뭟�NPq�l>J�a�ڈHx�f�����O�Ҋ4O�}�ի��g^���̤R��˲��؂,_'�>c��wʨ�J2?��$�Q��g@���|Պ)���$�Y��5AQ����+i�3{�E�D>��.L>�p��R'"�#"bm������Ř,Lf`g&Ζ�yʣ\�l��S�f�y[��웝��贱6�|j�?��x�mA.�";�9�M���E[Vz�{�e,�4u�}M/D����;�yXa���6�5*d+Η�am~E�t��Ĩ|$]	Pкٕ���SMDc秢�l��K= �i�.(�x�����PSI~�/*p'���kRφ(�����D2
j�U���/�^9ϴ�#I��Z�J����Tk4��n[���wJ� �`�43gs��B�?t9c�`є#��k��.��:��z.���p1�H*��غw�v��P�&���b�NZjă�e�r,B��~�䤌��3��"�k೏iv������w�JDg|�#�*\�H;*�eY�b5�t�f�'�ɨ}+-w��GM���i�:ڶy����O��q��~#��QF�X�J�%L�V�"��d��I]�Av��gh~��a��*u�>�Up,��l�͂B�:��6&�=_�]#����f7&B�llܷg{������E�m)C�����]�p��i��]D�/&1���nH�f�p�#�NCF�Ĉ��C�E��	C��H����V:��A��Դd�����9��Sf(��+�������X=�Wv:��77y9K3���l1�����:M_ Z��k(�wd�+z1н�#B�� �u�*��E�F ˷r���5��9������~��C)�`�J���=uѬ��DC��;�:�F�,�7��G&N�#�`�
V�̆��[d����zdW)���8_��"�sȧ�k�s*�+�E����}���2w��/�{d�� <�87�+ڣß�7[�@�6�iXKZ���_�V��;��!SX���P7
�g�R,54�����Ӝm,J��_���]��8U�u_g�1�"@\=��K�y�n���6��4St��O�@����ef�H�g�O�`w����Sm>w:W[�%D�8�΂�������F������B#p:�|�����&IԆUe�fA$q�m�T�d5){�!hى��7�N�*+�!<�.��|�qB4h�X�g��$?�=�pީ᫼��Q�v]Q��	��EBS6J���
�	�]��_�ޜ�9٘���������u�e��SD��?O�h6�Md�P�rs(J4���`-�iԝkX4z?����j�EП�_)bF�N,�$i��x#��x�����M��-��0�0u�m�E^.R�WK���v4CP�b�ùp�R�/?2��^Q�O�r�Y�/1�7�T��I�}ّ}b��8 �a ���Wa�0�?Q9�{���I��1���#���嫃�A��bAŮ���@z7sef{�i�`뛿)��s�~mUSY֗3��[�:�'��q�Yw�e8�"��hNLD@�����A�+2vl��VQ�=�ǃ;׎Ƴ"&�v}�`�����r	��Y{���:e�xM6yN=��I��Ɋ�	8�%��
j>-��틫z��N��d�K4����(T�7 o8�5�E��4OO<g��d'�rw�sݫ��`$G��,�Z��=���1>�ܶ��t�������;��S��*^�����&�x�J
n�\�s㚠�������tj��'�'/#�j	w�yF�B(ܳ�S��Qp���O���z)��{�%��gaWz_�0@�n�3	��-��5�PjƦ5k�v~�M�0�m��h �ǌ�B��Z<E/�Dil��+;C��*�7o�0��C���V�I�)�DZt�L�Z3�1��G�"(�[WQg�5Q"n)�K�#s�ݺ�
�K	�t�.���xѮ��N���(.rq,r~ql�#,Do9y�(�R	k���-����������T® }n��J�r��#���_�*��jF���=FsͰ��� ���-�uij14RM��i5Y�t�P�h;_�����o�.�m#�9ń��U����n�<?�c��J�R�]R.�4$S��P�����X��T��E�H-��ւ�,�h��]����( �߻��_)�\�`��������&��u˛��/eՅ�fSp����q�Pm4���ßK݌,>T>��;��12������g�>T� �.�o�0SK6��|���>z�ǭV����J���'��2;`4����p����7I1��9Lx����V��Z&�#���oK<E`hGN���?|����X�j�s?3]P;��T��c�C��>7�n��t/�©1F�U�\7�=�c�,���%L'%��u�v���[4�5ZW��s*��Fg�)���
8�g�X�`~�p�ɂ�tivU�?��.���Ů�[jz��:E�C��WNIt4�/��S�<E�V ������oWs:�"0��ʨ�!6;����{z�O���gW1��9�� ^Zҝ�����<��y��J,g��>�M��B��C8J|M�]��0��DZUb�uxZЇ�V�(ｅ��������J�Zѹ�/Z�u�!�{P�ux�!ue�K�����O�5�|�s�����|3��\kA�
��YR����� ػE|ZTXO��Q/}��"m�'���"�A�JxE� $�Z�X=?��Y^��xk�qt�a���Z��~��v�F�J/�H`{{��U�O������i�����+����6q�P?���⼩@ֲ����un�C��(9�3��B
̖d$�� 
�1�{t��(	�'�E'���cC�5k<wh�����o�X.z������{;x�7�Y���VWW3���W�a 	1;� |ﵓ Tɓ�u���z(AE����Uk�Scv��H�t��{q�ԍ�O��aE�&�w8����^�
@��\�2�u/T��_.!sD����Y��F�6;佻P���Q�R�0����su�p�K���<n�:����ذ�����������ꂴ	{�2Bg#�"�܄��5x����C�J:e-\�N\p" �p�(YeM� �b \�E��p��HБ4�r!�[�uW`�	��(�VΆ췇��� �ưs��(�U��e� ,�m��,m�N0ڃ��L�fOu��3��'򇢓��B�(4�4��k�ܸ
�AϬ����r[��I��C[n�%[���\����z_�W#}�^�^���cMl�/�Fe�h�J��э�ܱ�@#�ӧ�
��.�;���K9�#Y��@0�_�*���y_+7��Z�N<�֎!o({���ϧ}C ��l
�:���Y��;�rӂ���*�-�AmKH�㰗�D
%x5!�ȦA��lm~r���G�TJwi��
\���Pq@	�bPc�:hGJ��B���j=��8br����K�$�b�-����$��6������P3h+5�t
�U:�	�W�:Y|[�
U�j&������4�����1f�&z%�L����h'�#%6��^�檣0�&tMs��(��$�⺞�ks�n�>ϫ.4K��rPYR�8^�?$����rF��K_Z�8"x�d�4u�~Z�4�ƌ(��S3M0�ߌ�V)Z�>tWD)r6J5qY}�9��)(���B�V�\��`�=���^���aϝ37��2��X�IőAJj���LfRPu!�b�M��Ø��Bm`[V�x{����P&r��}�ع�(#�4�w���Z+k;{2v�&����LC��F�TRյ�L0=�IK�z/�dɫ��P�0�n�B�*4���g"��������{�<ؠ�N�=�
�������`�G�E�.�q�<zq&[@
vMFeÙ)�߆4��g�z��{��3���I=Z���C�:!k���k	�-��1�Q��I?�r[����,����{h�u�)4k��t�\���Y:&LA��Q��#�9��l�!Ė#��.��.�����薁��������:��ź���<��m�م��8�8��y�X�(�^8� J�BQX(�9�*���j!mΰ�]����}��s�)��7�\Z�G��9�2�;�b[sYd>q콴���c���|]�B����Z4��	���f1�,��0�[�N��	M�(�Y���Tٓ�q~~��A�W�K�"l�&��R��?\^����w���X��Ǡ�9 ��P��
��B���x��p�;�G��J��3����<�}����Ҧy�#�q�F�}��V�j�!�v�_��u� ��?�=˶_h��P;��k���}��{?��\��N����Mr��sZ�wLr6������f7�9����>��`%��=����>�!�AaG���O#�����v�I���""�����^o
.'Lx��P����D���Թ��Q5�$ٽ&�N�O�_�tw�����J#g�I��b$ƬUs�Z2^��1�~z����~�r1��.�X	�U�خ�}z �6r}�\��I�Y4Й��R+#�D�7�����Id��+�@L�u�����*W��9#��}�:Gl�@�8C��X�|� ��fx��*΄�4�lMx*l�q�%����?�M���~h7�&ד ��r��\�|�`������,�O�ٷ �V��
������0�w�s@�Dmd:G�sQ���C9���G�wt�Ã,��4IDE���!b���AN�V�* ��ɤ���,6�	�_�CR��:�,���N��:}�K��B���[vMFc��p���+v�3�����Y6Сga�af|�Sx*�!���U7�Te�����*X�H�k�򺎿�_��٪b.�;�������309��f~P�yjO�"<T���x���F��wtqB���Y���n',n\���s(/�i9���0EG�1~�B�gM�`w�e����j�s��\��ZOl	c��f�lrn,���>,� ��[��E̡J���R����s��S�1��Q��	��D�lZ�+S�dS��D??ؐ��̀�|f�,`��b��]:��V`���g��d�U��;��v�;���pM��v�����#S�R]+2�����,)�����zl�'+ �\k�^�?�X�2�[
����XvWl�?��|p���L"�w�I�����Ύ�p�،��@?$��ڋY]5���q��~����ܳ��j���:1rW`%���~��t��L��ua_�/�����
G�-/�@0�1���z�v�4�PŨ�q?%#Tm	���eY���<��c��e�_�X��^��A�F�D����� R� '7~��4p}��k�a��G߇� ����+;	0����.M�i��o#o�i߮\�"@�����y
Op�����֌2�i	w(�4D��7a1v1�	�>���ݞ#��V9>�u�Y�ӄm`K܂�Ⱦ>-��N�1�.�$��p�fL|�Ы����J��A�]CL�z�ҫ���0o���sy_�;�z�=F�W*<�z#�G lǉrl�_�D�̧������`P����p���+�U��y!\\K�/,�R�?�h����,Ǻ�o���2R5ܧ��+5ڬ#G���1�L���t�VUV{L�e�i�P@`�k+�}j�����1�D���{�7�=R��M��_k�LS�8��AI�f�Qs�	�5�zՊ��u����/��i�U�8ڟ��j/vY̘��Q�ՃuB��<�#���a&�٨�,��MREֶh>S������2h�Ek�6�Ԭr3���}�	*#K�4�Z���6[�����i>o���=T�r���͈�,��~��<6��J?�7�{G�y6����W aW�0~�����l2!�򦞏�+0���zt5a�,�q=!�'��7�Xuc�F��f��[%�
�$},��1),����-��������YXi�xui�����GK�̟�(�G��	��U"�~u��oF�y��>��Dl� (gBƒ�!��|����X�����ϻeN�{q������!]�˅9��h���!�� �NlF�Ipc�v3kw��}&�Jʖ,��(.:�TF��w������䕙���#�V�,�V���d�g�F��{`\rL�Ñ��fA#�2�u�ڞ����!Û�w���h����NO����M\��SkQ�`�t�ǖ��a�Š4�ġ����p��wd���_g��
��x��M�%J�9*C|ELdn']�ˊ�L�[Ŭc�� ��_h�`����Tz�b��Y�U�'�t���,��UQi�3Z��]\~Z�z!| F-ސw�;�7�&̩<9_6���/�i�_�~"�B���*Y���e�1_�-T�U��@��9:����'���n���&W��޲dn&q�n�TP�:"!.z����h�~�X�����5�H�?�`�D፱�\e~�)s��fo��9Ӣ6лWkN�;��
���= �m�O��͕آ��1e���:h8�*U�! 65��`Dbo�L)�Ar	��y��8����!O7�c-�md� ���(��Kg=�Q����!�Қ��1�����s����-�7gf�[�Ӕ�Ir���IĻ>�ݘgP}0h�'���3��H����#lٙCeg��%R�ﴟ$����o�I�*v`��O��r��q~�>�\%����±ͼ�q�˪So�]_Ě�V�r_��E�9d�(`&�n7j��D$��Εv����ۘ�����3��S�Jf�N�%~ݕ�{��ё�4��j��4����?�s<�� �'N����8�@;g ���՛�<���'��/
����5r�IS�_�E���oN�-�3������@���@��,7:tmw�a�4&}s����H5�ԅȟ���Y��B��eם3���h���%���a�".G�=�\�g�o8��8��"���u��Eb���&��LMw5���=d��I�ղ���|�Gd�W��N�w��"g�= ���aCls��w���$$�F�M.뿶]�������Y�%7�W���W���$�]�k�DU���{�fd�궲�X�X��r��
�IŢ�p�$� �{�c�����P�u	5]j�Q,c�/�cK��'&CĬ�^Pt��Z����F|~���"i�i'/󏗹4IL���s���ʥ��j��v�J`����W�/XR�J��b~����j}�b��9 N��u��/���WM��a�ߴ�4��%U<?0�/�ơ$D`k��}����2�.'��f��G�L���I���l]Zv΀�NJ����=�o�֢LX�}6��NL�G�0��r�Q�?>�M<9�H�K�Uۂ_� |�!� ���RS�y!�K��_�Ԥ��� ���h���N���q2�Ѝ*��������a�n*��7t�/]g�X�p�c0T��P_���$ʌ��jE|�4���I2yU�7Q��Z�V�m��Q�rɳ�^PŶ�k����xڟ����ډ�c z�'��(*4� ����t��˓�B)~���6�0�w\��X��}����P�] �{,�~�b�Iv�?:��r����^2q4�s��;-�#��Q��r��䕷��ف�+΂�� )�W����"L�����l�K��{���׉������^fթ~�Q�s��)��n�v�+��%��s1.���V�����$�h�E����?�W'F���f0o�Н2E�ʫ�uq��j~��R����#�d�b'}%�y2?�s�V�2�+L#@J>iC�Ġ���n��"��FQۈ�ؗ��z�(ˊ����,"Ѳ�Ueo�0�r)S�u��"|�X<kl=ϰ��#����d�@�՟+F��a���ۍ�\s�Fՠ��b�)?��_[��K(Ҿa@�]�@<K��>ANi�#1� ���Ut�i��g���jX����M���2��{ė�(�Ĩm˓Ir�PYg;=O��a_�l�m�y>EPkw�I`�^�^��dXE�Xf�Ke�R�y�B2��/ʪ?�R�����K�v��|��:u�]��=�����}�לZ�!ʗoY��%o� F�@!�Η7ԇ����K5��_/"�{�/�^� K!|��/x�f��l�t���A������[��&��PFp1�w�4}�;}oE��ȣz���1L��㞣3���ƋlMr�	��6�Å�%��&�D�Q���Kg�	wR���ݿ�E@�n���c`���3�� ���/��ܹ(.+2`P�E��H,�Er�b8��<Pt��w�����֪[�.݆�r���
���O��v��)��ͺβyǃӢ�Hf���;���|;��B�6$
4mj�R����^�`���ϻ�N6۟�i��T'1�n����N��A��9�C9P[��. �&#�rA�y�| ��`w�]&d����!`�B9nCK��w�S����x,�΁+Y��]N��$+NJ�6��J����)�ݧ3k�CƋ�N�n���xvƐx��0�>�x#����R��0�pc6ҟ�`��k��U��.���>��"$�[��S_�#M�Jfs%��"�6�̙�$���
�D�fhl~�(&Ipʾ=�r�Я�~�"M!���~֎;B*�^�
��>���=���^b��������	�)�7]ЙꔓdF�s�J��]w�ѧ%����5D���g	E�k�Aڌ��*G���Y���_Θ��|k������M�$�0�	+]A�(�m'L:B ���\�P�Q�V i���6���!8q��,,ѤA�N���3��*���)C��:hHt�q��J��܌�G�!%�Q�4�L�.p/$c�)FE<s&� ��Hgy59��7��P��Ct{�R��i�6ͷ��4��ˣd4��eǑshʈ�%�v`��BK�j �ڵ�wH6+�?٢��M���4�x��[\�X�{���4H��!� l��Y�G
�ٟ��B5[	�7#w���]���|CC���[��`9"l����m-
�K͗
�H�;
����^E����@�.s8]I]�?� i��K�~�wJ�6�M$���Q��])c8f:��\~�0b�m~���y����C�4�]���&�F��ЩC9(X�"A��%ҷ��Z��7d�VT���;{о1�:�MءU�X~B61���UP�Jx�f�%\P:dp�I*�	��9��=!D���Y|��<���s�����_~�&� �aÔ�$nHݔw��0q�hٔ�iO<.���v!^���h����kQ>�L���\������XrF�0���{5���̖\�r�8g nS�~���T�>]��3�M�Ad���Ddz���� ���̜�#F��Ef���:cj_�\0l�SBM:��]z����VHZx%O�����'��5 ]ō��'����U��]~��P1h��i1�=D�7#����
���Jټ-�����tY[�5��<_�`w5�b��Ⱌ�	}�B��ѓ������`޲���|���%f�͆��Sz*�/��,���;[o ��P��z��Ҭz���C��R��mzk�����/�5i�u@z+��B6�YW3�4�U�	2�
U��G2�G��I��S7#�4lfz�o�?E����Y���Y����".���Us�����F�"�����wm&=o���ND��SY `��/5��t�
�n�p!;}O.r�!r�9�$��+�i�?9�]9��M��|�B�����Vz��Y� �)��Y�T����k"MKbK%�e["#�4￯2"`3X�v�Ē�BC��S�ْ��\l@kD�)�kDdO�<�����y�~ѯ��N�}~|�H!P.�\iu�%��L��&^�v�Y�bH3���Wf�k���t���҉�k��{��&5j�������[?%�D�5~�j��85Rz�#�h���=�/�X7w��u�S�B�����[���T~�P����ǃ��`L}� �/J~9 ���4��F�C&��s�r%�:J��i�8�Lrq�,lѓ��Ĉ���U=�4��]7�&פ&>��T�`�X
J�$;Q�0C��߻�t��x�I)�`����Z�X�Ư����.���+ր�2@��b$>0K��:,7�/LЪ�u��?.u},Kx{�N���ܔR�����s��vߚ�s|=�b���}Y��::�p)���޳vP4`@�8$�<����0|�i���&���u��@��(v�N�B��:\�DmhW�V|�����1�pW���i��@��?�X���� ����aΟ.۵#v��+Xq�ꠙ@���B�� ��$4�����	j�K���~$H��ONj�̏vq�0�{���p}W�}��&ŠqP���I�W�<��佚n"۷�
O��o�I�Ձ��ށ���$��.RT1�4΅n�aa:T��`�d�9�մ:6�bK2�(~��ZsQg��A1�ú��afk��[A�\&�;0Yu�,	�;�	�a�êp����׿%���☉�&�Y2�Q�����u�l��U%���ʠv_!}N���g�)�~m�5��T��C��AR�,Ę�N<�)9����،�U�-0��чi��T���r��ֺ��e�A�:�=�>������cY�ۏW���^usz�iN��r��l��#�Uiy�"��� ^��.��>���c���ͦ���A��)�{ʂ��A<N����D���֑�3 �^�bUz6�2䫂�@qs����y�����/ *��#�[���)�D�=,!�E::����-%�����`�Xr��6�����A��8�ݯ�!+{ejC�x,��yEm�@I�>
��N,.�S�9��t��Pe؁>؊y�GF��Ns6c?� �{��gp +2�m�me4sY��9���_CP���3�~Թ?���g�-2�P�"��D�{���D�c�$+�p��p�MB��3��^�l������A'��ߍj8�t�F�I'���K��h����BB7�N���S=Ŵ�9�-w-�=�S��q.�|��J-�sy�Z=ܴ����>Ӳ����8K �[$u[RW�_@�a�_x���K(k"��W�� F�(U���9<�{��-L����li���~����G����_�V�o��I�uȍ�(7���hxg��S-G�*Z��TS��`*�[hxyw��gzx�P$������T���p�a���Jya�k}�f�d�y��=� Ʋsk����l|:��)v#&B�dI���g�ʋ��˝��(���K�d����$���*��/Y-|��5l�ײ5����@�2i��Q�ӎ1���VF�P����%!���@H�»A�����%�R}A�܊��r<*ZLj]���{��r�t���(N�H�<Y��[H�NQ�eb��lN�	7]^�~ԣ����	ZW$g`3�wHI��G}*�>�1�.���0�}��h��!��<��P��%?GH��1d��M��'ں�r��т�R�����Pz��\~)r ���/Ql��!��@�D�-XV>�,�O�-���T;_�a[q'�������zG�8����ʘ�5_�r���Nϝ^�R���-��߂mB��<���� ��ך�6H'�x��Z��5<�C��|7���Cp�T�bǦ\x,���x�Z��^E��L��w���r Ѐ@�"��Z�`D��JR��"�R�a���Zu�.��w[^�r~���Q:,U-.j�&�)��'���z@�֠�[?ds�>�N�^bU\~��U��{H�������D��%{����'-y�혳�M�L7�>.%�z����G��������jTs�m��9����u��=�b5.g���Y��	@)��̨ORp"#����O�����b� �Ь ��~ʑ�?���-	oR��u��|���4��S>vY記�r@�kcĄ���lX;7`��g��ֽ8ꢄ<��/GL�DU�h��Q�5�#�7�}^ý(�V�3U��R�*D�?�V�j1cǄ�3;���sI,��
���Cbrg ډ��S�N%�!�&cA��y�Oa�����S��p�#�ü�mg��M���R���q���5�͖��f�V%��i���&.�Ux�D2�e,0��.���������������%���� ���تd]�bH`���J/�)Cx����^�u��#�jϲD�ZpE��~��͓�ƹ��mlK)���+]�-/�,��pU���*1ב����lT�EV��Cp,l�时�%G�Q&Ԁ����)���+J"k�Oޥg/��Z��,��@]����U��g_ysB+���"#���d�ɻ�9�3%�6�dQu�h�xm&dK��	��6H�<�yk��U'1����{��(ci8`@Ϫ�K����6l�}*��MRh��`�!�|�F̐�r|��kE�Y'�k�����d-=0@�����ґ5���&�D���z�:�(���H�R>Rm�c'2�"ލ=f斌���R��+����3��_�კ[����'{��J�EQg�n����f -�AEÆĞF�t�)��"������R�i�E�z�� ������.�7��y1��֍w �Sh�a�Z�/�l�>�)����R��G7rt��}0�ۻzc^ņ�	x�����r�"v?i�k��w�D���v�NK�GrN_R:g-l����̄6pAN(-4�D�����
Ąx0���H�����VPs9������f���ޢ��R]ի]-<�`%n/�QL�hA)�=��������[i�i��laxs~��NL�_jMO�U�Ta�y�;�a�*V<�=�9�W�9o����EӐ<:=�o[Ch��-�az��'9e�f�S�GWf���>wnC&�?�bX8j�؍!��v�dZVD_[�

ʰ�Rw0�9��"`�f3b4�e��MV�Y{���pv𪣮L۽���3���X7{Y�X��̱���Q��Qؔ&�q�C���ѸW��α^��y(��i扞�'f�?C��\�h?X �UG��zh������X�������L]��Q�=�? 0�<�?s���c�E�}Xq��_^�+r��Px��7��%�y"�qC�z�aN�P㬔����F�M�OcZ���@"tdW�����M��Y{<���V��v�#Loy�KVw��!�:�?����L#�����|
�(�J��`ydf���<��q�&� c
��$��q�® �a��1�_���04���dɡ��3�Ձ/���?sN������[s�V�5��2rG ��2&�[���:�ֽ󍉋`jv�ZE�|�Yrs���F��	�l-�������]�8�o�a�F��To%m���F�mt�Tf$oSv<s�#Ǧ�;
w�+Ǡ���cC�ޠ���lb��ʼ[�S��������a 䂲�Xs3��܄���4/|.�'�A���j|�f�2�{c�o~��ϛ�ƈQ=��:&(4v����bD�*�iZ�[T1>�AS��ܮ]��.�@7&�w�Yo� ��QV�%���J��Cz^H�}a��ܔ��0�.�>#�!N$_���d]=�~��Η�R�Ts��~�\��XV	�l�'�UI;�!��7�u����'?��+ ����SOtb�'��HK���{����!�-N��@8��'��E�x�T��a�u��a�|9��b�#��!&N�q�|_&L6��(伸f*�P�z��(*��3��I����'\�dJ\�iVzM�&�K���~4러w�Sa~b7B��Qeㆦ����3�TJ�K�y�n�z48�.���\@�)h���CX~�q�d�CA��ko)hrwI��A-�F���*���J����/v�Kv������Ut��kˆvI�3�N1�3Ki�$��^��,��Ɇ[��E�0��<�xj�i�A�D���7ۙ�#��ь�{&�"�F�%�7�ϝ����+�
�a=@�*�+o7 ֪��[H��9u��"BAy`�����ܒkr�̡�� ^�P�[�4ՠ��H�n���M#1����j�x�����c��Ӧ��m��8s�	�Ux}vj��.0S8e�Bt�Ë�V���C�� F=��C�i9�����̺��y���PX'�f��&�p�Cn}�5�"���A����-mW!4 �� �i5X^��K3T��m~���.͙Y ��}K'XK��?܆���lV�_�,���� 2����3ŋ���m��2�]��%���J�Om��AD��Tp%���G==�p(qX�e-T��iϨU����3�i\�z��kdh��{&�1�x�S}�+z� �q��6�V�Juw�If�N��i�N��H�(@Q��vG��CsɈ��e�+#as��w����/%��#g%yf�:VSF�,z���~��y}������l'��P<���4��E$7&�MTIL�^�����@��2�O%6�0�5ڟ�VE�7|������Z�k�����i�',�[3��qv6��j�q�2��":K�+T��ڔ��D���#\����>��-����2Րݮ�qu���+PT��Vg��z���n]��1Z`�J�n�v�O<��3��������<�F�(_�S�d�(S�o����aCb�P�SV2;�2�T�K���q�KK1��̃G��s�}�&/��X݁�v����K'�d��� b-�>�(z������3���{���X�j��~���Eն�@����=l�M���>���;Y,�Њ�,����q~ɐ�ّ��ר�A}�"������g
�aEOa�y02��?I��
��7M]��Ȅ�4	�}ok�!�/���&t�����|�U^/��5ծ7v��VϮC+oҸ�J�M�l9����4|�>KU�O���+7�`5���8�}"�˂���a�3x��zt��-F��79$ʮ�������`�Gd{��@A:f�*I����>D���� yt����j���	C
�3K��L	�`rԺ��͕Z��ڴ���B2G�W�S������ԼT�YUwA~���XP��'�U��bA�.O�}�&O7��y�)�7c�T����kn��H��=����Y}������Pm�@����W̽"��r3*Z޻��ͥ�	��K�q�ﹼz�|����p񀬑ݝ7^��K�J����L�:vs[m|��ܓ8�p$]vR�];��p,q���m�g�H�hX	�-\$Յ��L`
Ccƒ�}ym~؎��=?lT�qRj��5��"�"�G7/;]̻�K�k���qp��M�9�>=/�n<���0x�)�x��L�-����b�MX�j՚2��;Y�3򤢁�.��(���~��0Y�C`3��ʺ���+X��D�}15W��&b�8��]��q+S�3�� w�"�b��͔�a ���x�öS�Z����������g
�P ">0Fvv��`�L����3�`��G�q4`y��m �.[�&f�1�k���v:���y�:����E*�ܾ>������S��Flm$T5�z�S#B����>�O���Es�kn~nx&�5� %�� i�D�T�׉�m)+�\~uNb�������H���"^~H]}��]�O�i��@���5��lwa/Kޕ��}]X�^�!�+k՝�D�9���c�_�q[f�  dZ=�͇aHLc#A
޲�P��{�
�L��1ְ��k%g���R�(�V�s�:�P�(�~Š�������؟f>�������C�Vfo��Z=��?��D��2��B;��A�,����R��6���h��bB����i���ae�]@��� �J���N�����@)��L
�ۉL�6�^T��r�@�5N�+A,�M�6�S�*��Da�x�l�Z����|ԥe�~� ���h�9��~1�|W��8Ww�/z�@�+|�]v���o(y��w�}�m	sɅ��#过�����ee�ci�����Ә�`
D*�9�'�A�m.�~W<)�{�{#�T���zs8�;\��f�,h��n;��,���d>�ܰ^]R�� _� ��{��yUXop:�1��+]�f6���K��_I"2TS�>���b�e��'�E��!�V=a��>�e+���H����G���}Z�DU7�;�0��'y؏3sZ?|�|wy��J�hbb���(��/��8e�<cBM:H^�Q���������7��0'�.z��b����tͯÆ���F���QQz��C�+ ������R4#b�记#t��W�'	�^�f"��q�
Z�a��>ߡ�G5\]���x$"��UP.����0ϥ��٦���G�[H��e=�*kN����nHAȳ�rފ���y�fM_m����m�Ϙ��	2�P�=|���(Y�In܇U�p�%���Y�T�S����Pn>!\g:yc����b���Z�u��ڮ���5��mFe�H�k$qo^[��X�5�x��tm��Qy^@�������IW����������f"�<��SI�ߒ��Z�03N��8�zֿ� ��j�%DG�F��o���s���L��2��HV�����d3t�x�',������UgX'�r:���:�*��fU�A������EG�X���(�A�7!�Ֆ琝P�|�V�p�
�5Iv��;@l��qAb-��pi���%���@�ݭ.�r�=�w~T��f�q
6'��0��U�� Jq����G2�d��M���Ɣ}[L�Ӕ�e64}6k�O!C%�.%U��3k��<��g���\�9��HB$���$-�G�I�&��1%)�����~[�����;4z�����������ܞ��ϽJn���=a�9&�O?�뮠e�H:rb;�dB ��G���({"���\�L�.���V���Q��������lr}V�r*�.Al� ćU{�zwT��+%�/m��-�� ��x�)o+�U�s�y��{}~������<��,}ʧ'Ն7�4���+�����ڭ��5�^k��So�N|��]mfќ��Xw�c�5�my���h�<9��C҉��;;̠Y��$����������dc��M*���r:�TS�c�8��#)�dt��H3�̼�/2�<�e�~��`�(���Y�����葖&��,
�͙~J~��T��Ȑ�v�b��<l"��Rm�x�ښ?4@���<p5�����7�q�ДH��OM���$rI���DC<�x���\���0,��'�@[�����f+��1�9'!(YQ&iB���Ah�:A�n�<?Q�IW������g��ņ�8���> nXTM���z	,�+��� y}8!�6[V{ɟmZ�}��I�	+��$���~^{�t�N� |����u�Q�c���r������� )��6ǹ�}z�08Cx��4x�|�ĩA ��&]�d>=�g'2�Љ�)e#�X�>�0Һ�T�v�vT��;��V�àt�h��$�ss�i~� +	A`%�:B���E^��,���s�t���.�8S4��������+Cu�{����VЎG�!��n�x���nXW��I��$�E�i����+e�"����zI@$B�&�_b�N�s�}�U���o�E��^,u�e�ɝ�RPD5
�K�n�v�AX�ʘ���D2"��0ߩ��#���s�� vp-I(|��.^���b��E�囍���P�yg�C��մZ�h� �9J��]*�?d>^x�vG���Ǐh�hne���1u a�p��l�]�6>*� x����S�jP�����W���Bc�96n�v�c�s���3o��x�aLo�Ņ$� \�2�k_��@f�:��#zhM�-�o/�4��}_	����X4�Hk�_���4D��A�t[ ?I?C�-�c&���A�N�2�����P��ǣ�vWW�ғ����k9N���c�d��
א���0V	E0 ��������0�a��˺�i猘�_�j,�cfxV��WUf��a2�l5�*ه��	ӆy�	1��)o��'6�f�Q�����5�g��!�ND��q����{���H��Q��8F�XJ�-�>HsUB�~�I벳-S�����_���h<�
}cM���!���HO;p �3kW��@�\�$�J-	#.�:�P�2���@���(�MI��,9jY��Rpe�|�o'�a��mY[M���*c�NWN6��R����f�?K�Y�\����,���c�mH��E��q�~��T���F(R}Ӽ.��)N_̟IN)C7H��Mѐr���6���T7	U*��E�_xבl�'.���ِ2�4*N����-0���jw�F�/(��PC�/��]7�S��h�Yfۃ����]�Q7�$M����˲�;\(tYD�%��e��1�< ��pYZ�}�,8os�鯦9�����}CG��uׁߏ���R/�1Kc�7�����N��z,X������gE��զ��V)j�� 
��e�Q��D�-MK��1��ؐ�{�rUa��8�tm�j�;Za�*����������Lkz#Č�.[���v��MU�;4iEP�:����M,"�d ^�,�9�S@$��m_���5}M	��
��8L/�u^"¤�e�^��ܥ�ح��5��z\V �\R�U���T��H�o�\��-��!E]�'&�S�s��cz	��Xi�W�yΫ)b�(K��9�u�a�'�*hW������+�����^��41W�� �k�����s��Yg2�����*l�f��pG'e�DTi�чޛ�s7�Yf����OfG���Аw�%�����D6�EŻ^�eu�K0�b���@,�1�H'zIjR�R&��dM
TT��2$'����G�V�}d���r
�7s���xS�auA��S	��N��ړC��R0M71L=&�����Zj	;�4Q��[��~�������s���̭���y2<s�s^doW���"nT����V1э�d�W7�
�-�cQ��o�jm�i��1hap�u~�s�B��!�"��ٯ9� p�6%�Nbt���)-S����X]i�X4wg�������[fbĺ+H��ӹ�)��`=Ӳ�zh
�yO���)�� �l`�����a��T�52�����d��v��J�߭���Ҕa"6�֕��'Mi�'x񤰑�>Z7�K5%;[{SG��[)�y*��^�df$5�����װ�*z'ؽXe��&-��>��9  �~��Y
��}h�a�4����o�>�H��DB���Y�v�`��$�o6�$=�3�Vɕ�&�~D�z��4��m*�W3ܸ��HQK�/�?���y����a���/,�u�Ď�3��gηK1��X�r��BM�p��m$�ˤ��K�a��4t	�ji�
�u~J�e�fv�%n!��t��8ߏ�_N�`������^x'p�_�r
|g��O�	F��~��&iWWS×**�+%TǛ_���s>��aL�����.y7�\��{1hP~�!�����|����z�`�D#nut��4��x� �Z��M#���~�H9,�g�0z6�S���n�����q΍�CHI)�!��P3O��̨�͍�(?��e �k+�}��!(�i�la�]>�`\(k���U�`Ը:/�u�7�T�h5�f��0�p��t@��GuW�}n%����^�j.��w�v-�eS��8RC"o���"njU����|l|)x�Y��r�CD����N���/0�O���eM~LM۰�Ƴ�A��uOJO`��?K�0��S~\�7���,��#�g�;�d��F�(��ލ��IC��m#^//��W���l��p|q�lp�^d(e�[�����7 a�0[�-����Y�T�]�0�dyPc%<�.�c��K�?ͨ���$!dG�Yh)F��
f�3��~H���
�x|�q���l��n@ޠ[�=���2R�Y^%;�I�Z�^?�C��j�RV��v��)��ؾ���TwW;`���+Ҟ��6�-1�orAm�]VG���*�?��-�J��瀃��iR�lvőpp���\R����R��?�F~S��[1:�,2�Oi�"��]>b窺
	���4��c��5��&6Xք�t��E���U���W,��?�'J�	�{�tM+�s�Vl������ֳ0n� � ļZ� Wzz^)���u�Sr<�ו�8f�-���-x����� R�s��lV����eF�9& j8|�6�����l	^�� m e#�飽	_���k����%�y��Y�x �����B٠M`S�O�k]sPo6X�hx�{V��r8��L��.���J�l�.��X֢�^���^�� z4DtR�	@w-3�������,˄$��A�q&W�DC���~b�ό���79�}�ĻH�U��ښ�,��[pRy���j"�������`�����6ޙ���mr��nI��_���ytk����4�]�k�G��uq&��.�r d#`�
����M�fD��^����t��9g����X��Gx1<�3�yw����L6��Z
b*�]�L�	f����)+�\��q}VD�w�;�]5�s�C�P�2D����A:�͵��:�xR�ȁ�Z�O-����yš�9�*���V}*Gp���[2�?�U�gp��J	�;7*>j�$?�,��(><_����A�F�H���4�՚�Q<�0tI���(�||h;��(���Z�v� �g��UO!��F�L
������7�t�f�ʦ��`��mQڹ���*mL���P�`j_�Ҝ����n ζR�-д/Z�<FN�v�����ǯ��+�=����z��ef3�6;Q�GW�V�G񱠸[D��ݨZ7��L9 \xz���Z��������3E��܇E#�ǳ�DZ+�rXҏ�N�v=oH��ny�/�O{��KuA���Q���4��e�̋ ���*�O��2Q�/Ϯ-c��=�/��)=�^�ĝm���Ž�E�XH�bu9K<����5��D���τ�t�����r���I]kTڮ��ل��U��V���[���O-}�Q�3�cDM�YQ�_$$~��J�>�GcjNO"5�Q�y�&}V�-F�l(���* zĐ�l�ŏ/k.���U_ �4�p���D�����ؿ����ÀD�ĺ+Ȍ��Ɂ�h�^:x��J�iy܂�����=`��W�p5eεO�~:������ �1�<E`�H�E�&:hHp�:y�� i�+$D0LO��0��\T��?g@�;�/*v_p�(j9v�u_��ߴRj�
-\�~����u������J��.���hzd�[���$�������N?̽=`�;�\ �`�V��}���jֺ%��:\|�G�‎T��k�[��xp�a�~��d�S�s�X�7
�����v{0�鸪���k��$g&r=� �:�z �~/P�S��&�#}[DPw��J�_��u9�/jaD�me��9j�t�R�^}���8vQ�Y�{�ۮJZ	nE�7�|ta<1:�\��Й��J�i]�2j�Ui�j�q��w�]�����gb�(8	N�S��=��$�e%�7'π�!�v,���]� �Q�������{����J�n���[��p���������3=���W�o�S�^�\,QK��*��n���e���q�A)Y#�S%�B��]Opl-$�nƁ��
]h͗B����_A=�_\���݃�����[��fd��`������L��aG����]:>�amg�Ab
�	�]�Gp�z����,��`�o�ی.-�3��`��S����B!%�ӞJ�s[IGޛ��KhW7�Zp��������9E@n���s�J ��6ջaے�����6,s�������߫ܝ��uY��ٍ/y�1�D�"eign�WrH����A>;�r;1�{���1:J�SEɞ��[!�TP��2�ϛ�)�Ps�P�P5I���T;�抏�u*�v�.��&���pj���'2��Aa��^e v�4���a����Ϧ��l,������7MN�-�����#V��H/�F�~S����E9-G�Z���Mn�?k����Sh�C)2�t���'k=<*��������&D�=�F����r��1��m��̆��d���ϐ��އ���rB�:��*�d�FBL���7��˓�"���f���d3*�)\l~X���'k��^��c"���a!�y��%�Ǵ��=��&�Ɠ�3�:�����Vf]�_!V6S��7�9� ������,	Ƭ��v�F�Y��tsn�6d���G�Lp��n�U��Ho����~Ϟ7>��b��y�pN-&�����F<*;_��D�v�J&�`��� ���D� �cgeHa}��L�7��4����C�Ǒ���n����F��k���=,;s�&.I�|��+e����SX���%]������2�y����ǩ�#C��ƙp#eֶx�vl;j��h����Ȧr] e�(|�?Z��%�T��Vm7\�F��+K�}����щ�кx�
�Z	�#iz"�iXг���F��؊�
͸�g���Qr���d��Muش�6O[uK-п����}P���!�\f �n��Е�q2R�0kW>��n=M}��"|���IvB��3PC��5�d�,!�뵯V���~Z.�t!^z%���I�b\�v�UGwU�K����/��!L��˓�8���V�Y@g[4�)Q�r	��fX���I��hSyE�.n�-�/��9QO�J�Hm�k���т��͹_��x̜p�����+|E0�� �ǃ��!�@S�@PX�h�H6���N��p����b5����e]@��8�$5I:�]� �UKd|~g��v�1���67t0|UA�2�6���\`4�G+t(AE���������(Jx�wFd�$t�X	��CRvhD#�O�B��?�q����V��� tt�Tv��^y�=��"j�o�L7�0�� =�=Qg�
$x�ҳ6�F�~��F,08�q s��D���;� X�Ϫ��m�@(�o�F��z���d�%F��wɠ�-��sQ�,ʷDMGOt�o[�_K�ҟ�kt�R��ӕO@rx��ǃ�����v6�=��s� �  �g���Ke!�TUloVO�\~8�����}���۵y◝ؕ�A�Y��8��&�^ʉ$�n�;yМ�y�j?H]�Ғ#�`=��sӈjyY�ߩ�E�DO������P/T��a.��g��W�ʌн�˱��2�-�c���y�|�/���[��7�y�yt7�T��^�����O�&]�r�	!A����W_�EL�N_�
-��٢_m�S��4w�؞�[x�d�'�NT6VPk��j�aW2��MQ��nɉ.�]�sۚ�I�ӹ�"��6���x��yX�\IgZ ���;����yڞ d���L_�cY���b��p��ȒsN��8qT�Fn��pR��Gp7'�(�l����S�|	+?#̢D_O�818�}�c����O��P��Pz1���$������!q�w:�x4E�Sq�o��d�~����_��7�k� �U�9@��������g�h�9�>�ᴹC�'���`��:�ґ� ��k�|{����?��ݟD`"��8�$��N�V��U+:�nzSc���vD�^h��KcX߇�偙�Y�Kv¥A~4����=������OP���fŬ ��M���I}�b�*�)$l�<�[���p��S�����L�M��[��ܛ+��z�,[�'wd�Y�hbt�f�yK]���d&)��42_���q}�v��ܐV����A|i�
���Wr�����F���tK�ka�D�~^��q���ڼt�N�>�݇L�ku�`���m��0U��d���U�jq��c��!�� y��N�F%n,��2`����Ջ����'��L�Un&'��Ú1�7*ȜX�����	OM����t�T�W���� ��r:b�(kaJ��������/�yo�7��÷�mvZXѢ�>葉CC�����S��26�5^)ݏ۽���Un�8ҼX�`���0;��	�å�@����뮝��5Y�&���3�Ր��/��*���o�U)
]/��VE���`�r�-;�Hm�.H[�m�H^�d���$_��9,�Dl�?K^��D����S��"^��P�zb�Tw����z��')<�>M��G�l�S�g��y��?K���md��-I����a�p^��@i�z���n�V(b��x�?}τ@L��,��`��) �F��M^�S��D��Az������uj���|�4�_���I����ԮT�����(2�xn�RHy�\4x��I��/Dre\�@��&� �L�m�BQTe�fw�[[5EE=�A	�k(���&�	�L�EաBY�)6��73�L��$�#�l�:�<'Wt�Ì�1�����P����e3$���*$�6{��Cl���N�&�q���Ħ*n7��.f-/$\f2m�ʧt��Ib�"2b��B��o��`}��Ӿ�j^�뽏��eP�#�ut7A��ϢGٲ���/?5� #){�È��]xg>�J.0�����űNNt��8-���⠄ך���RG��/-�Ë �rnoj�"ѱ��m�-3j_�&ݾ`�UCY�k�j��
R��n"�-2��7��54�O�r�I@�
2����5���|��ҝbCe�F	~��G���2��x�y
�&�^\ɾ�U]01��S���h���D+A��G��|3,*l����+c����N�}I9]��bm�Yߙ>Xu��pۄ&��V�s�o�{�>��`:B����U+F��c�Lޜ���yb�@���
�p��u|یX�G]��`d�Y��H:����J��ZFV���'�):��e	�*��J��Vh��/^����v�M�K��\Qs��-��?s��Ar�u����ȳM,#-���C��h?r�~�p�9�l�ͧ�p0Hz�*���a��/�;���h��.oځ�� ���9��1���ڰ�> ���8E��?�������Xxݜ~1/P�� ��C3��q5K�cbh\�f�Vx�!aB��r�g���9`�~#qݛ �eb��d
��[̐BVFt#�Ͼp� ��8w�274���Y��P�Oc��߫��p���-����Jo��ef9մ�������,����z�a������m�u���)��#�Ky�w����*t#N/gD�ܶ��Ʋޟg����{��?�� D�ބ�lI���+p�q�^���;87h�"`fOc������ޗ���6[�"w��3X�uЋ��T����Sٌ/���	��+���*Q�A|�9�'Z���K�jM����c1��ʾC����������%��I��@��V�]'���^
28hѣ�*�:n	�0��kl�>&s֯��-t�q߅ҹ����+�˘���A%���%M�o8-�ۏ�.�M���xJׁ��zh�w�U��BI���x	����r�,o�yv���`�Z�i�ۥW_Py�u?���j��J���]Gj��z�q�K|��=:Iŷ�H
�>��WN��]L-�P�
!퀽Y�BK��85�w����&��]��%�9Wէ�H�����b��,C�KB��>�;�惭�j3��O�g�^��(|0�o�!��e����\ѿhV�g��a�9���������p� C��P�P�6+{�#Z��H?a
�b�`Nt�m�k�����.��b��"H��`�i'�]�y~f��B���l�����܋/������m1�O@	.��V��1��3�eM�;�����b�	�0���į�T�1�"�c�z���|�.[ #QI��w��b[� j@s[�x		d�ɕ�@#�6)�ت��T���%e��0���Ջf�&� �8�i,����L���W/s�NW��&X����/{��S���#��Ib��R�t�4еD�B�VO���[�U�أ���?Z;�����mA���|mܖ����K�>�#O�����k��������),�����{!���@���Mo#�����Cᰝ�-~i�{�a;�kɖ�� �VJ�R&������MZr�ş���>�u�H�ĉ<O��9]��ݍ���DL�dfw`#P�R�y=x��2�-��I ^�����=���ҋ`��'N ��B}�r�ʢ�y3���*��~4p��t}{�<;�y}��S<�qAPN�/QM�o���;%f�����E���4D[G{��\kbϛ��n��bkN�����Q��b�'���<��R� /1������C]T�1=�n-�?��S�i�E����]V�ftr�����:aO���d�o�����aѣp���h����qS`��-"�O�"�����R�����x��D�1ۨ����g+���Q��e�����j���1�v<�p��o���|�0�8kVw�VU���*�=h1`�n�_�m�|���-��&6�Q�xX?��-Y3f����A����>*���U�}� E���-@�8#_m <�h� �sh^�)6 ��M;6�7�"��A=�lI�$��ҁ�,*��SPku4�hiz ��+w~<�ߚ���G�h}���F���O8.d&������%�QvF�9+��D!��z��n5�3 �~*1�e~k@�ez���\�*P�{ԓ�f�R��+�%R�o�>�R�T>��,G:'Sյ��clZT�6�'���Ss%����b�I+E��n�
T7g���2�	Tf�0{u`��N�=��g��iB���&�y_�G�+���&��C�/p`���gzQ���ieO�HɆO�I�	"hx*f�����de�~~���d�e4ب(����N%"]��A�_����
/�>%�{�ZL�"�}��?s]-"�f���B �(���c���m�MS�4��f���FW�99)iDx���x��}����R�H3��1���0�X��-��mV�.�v��><�N5�����2��ܙZ�Ϛ�;���#���넌�D�\�dé�����Q�ю�,҇>���٥+@6I9K&��gQcFT�T�b�yy�(M\Ǭ3�xљ��J}@HK���a�Z#�$��#eO�n'�	%щ8����%㪦�Rh��n��K(,^� _�t3n���y}<G�a
��+��E����<�2=Gw!	�`�c2fLۈ�g�c����mG⯮���8�V��Ϝ�ں�5K�p��6���Y��ͭ'�2[m��Co��-$Ϟe��}��~(6��ZdIV��@����'I�P�$7�v��:�h�h9$/eC�����D���wm"S������9�+�6�<�[v"p��S �Cy4����U~ߴF���)�$���K��� �kz����1�;|#���'db���:O�ԕAAŵL��j\�ӳ2�^Z�e� Br�pY6؃��E�.E��{�U�i�}O�4I?�ʹV�kgE�8(�v}1�&��6�3%�ZNR:��X#�=���!���󈖚��&R֌�P;3����F�'�n�"!��[M��[�R*���}��Q@1����zk���-�te8�!��@Cs�5W��j��K�~<�ߐL������Ԁ�ŋh%ċ�9��pz�}�<�O��Gs��Qw%u.��%E��1�vn��=�s���FL�|�?%�׫n��9���5�3�3/B��I�;G����X�?X%���jɪ���9�A!��IX�e#ݗ�p��q���W�!!��P�	��
s�E���i�萻<b�̠&� tYʏQ��;��!����g�i�;d5�ەn �Q@�=>o�����-�kF�Cv�@�g��O�b6�M��wG������vw$NP_��_�
�� Ð�brE�9t��_u̡��`��.�_�L ��B�j_�f����pT��q�-�QN,)Y֨���p��l5_����{V��CJqZ��V�vP�dF� �o~V���jIpK´��wa!�-��aڧ�J����oo(j} �_I�B���������*)b�m�+_>�I��~���8%�y�%�T��E�{�������ʹg�������*�N���a�����ߙ�/DB�bl�+'3�Q�0J��Z�d��%�/b���3�%E>�6�{:��2�ʎn�HP�O̘ɋ<o����/'p�����_u��t2��0��
�"�Fd��N����)9�)��TC��_-JF���W������_����诙	�z/w����g\[P̾�����l�h
�Ђ��6		�6��U|���`����h��>�Ԃv�Yl��k�q���a�U�D�PH��Q��,�_�I��Pz��:�H>�O��������`�M&k�jډj��ZM:�\�xlV���l���2as���}��k���ղ&@�V6gQ?��+�kI��f�,hN]�۸�X��^��7�c��]�[��
��|�g")�Q�Z�NYTʔ$=�4�g�hہ<4��adI��LW2��,�����6̹��fF��,���V?�\@���q�glbx�Գi+�b}/6RY�Δ
|�����Oi��,b��A��@�BP(�:0(;�3�y��!�<>&�mm���p����V��S��m�Y0Z�m�ǉ���j��E[j|�:4Z�Vߗ�_�Ek2���7�ѵ���4�"7.���z��&!~ڛ�&�/KAW���h�7b���P�C�$�aa�t�����Pu��P�z]��C��?�:zQ��{��]�K�	� mtX[�����\/�|�����&�J8��}hF�$��!~ǻL*��*�T�B�Y�b����'�̂��2��-����s[]��Rbp:)b�#�E���AH�U=FU�����Q��(J@p��B���Rq�se�E�pw�S�Rn��as�P����!:J�))��W�L���hT�<P���������-N� 8l��S̏FI���TT,2�d�i��'3�Xϸ�H(f���q��i*�}��Nh�?�ַ������Y7 _�#�}_����m��e��V���e�S���?�}���=�O��^b�9"�nK��V�+�J%`:�6\'M�Z�}�}>�H��K}��_�=e���?L��3r(��/Aj�DN�=��Ps��J�.�~F'�G'�yϙ��acS��-��g�B�	Ȩ��0�]ɧ�B��ƌ��ά�'~��D�������Y�Y=��8J�q��+��"i�{ <��\������Xh�������j�m�[@#U�_bZK�?�:��Y�'�A�e���O��0��3�������(�:�	�g(�����e�#9�\p��.�_"gK��7Z�c�7괊j�EK=��!���1����`[?��C�]��~�����
*�\�3ZU�f�^��	F$�>K�'�g��	��T���o��!Ǯ��Uw�\� E�$$#-�=���ܱ=��:�J��C��"o��ލy���U���������<��	��F*{��!�_�Bi���8Ic!0�{.�$y�7w�ޒ'�g�;��,�d��CW%ɱvYLʕ�B�w��#�K������SPoǻy�g*����3�c�pX+���R7������.��&�����# `$
&�bV'h�-zA���E��i4=�wl��g`������7C�l�ޒ��Bϗ����0-'��2��K+� �s�9����Wa4x����{�����"����&�V��T+��VǽXQͬ�Z�<B���ȿ,��K��5�@�~~�č�Q�a�}�R>���Y*t���D�1�]��ݮX�K�A�(��/q��<�]a�|��Ϙ��p�b�51%���0���	�U͞�;��pQ��h��&A���ҷ�B���������^HV��o��<��]f��(DYE���^�*����t��6�vhc��-F����T2���N-�!�S����+��G��n��S����I��[#�{���[��yyES"2�=���1裱���w���o)�s�ń�g��h�Xd�q��)�P��/*SP2����U�����C�e�w�'0[1��7H�-ݮ]��*�������O'PK��-�eu��)����}_"�S5;@�,c{�V�?+���M��˼n�����
>�%N"_�K�V�s�"���OH�q�Ԕ�g� ��$V���;�ީ��:��)�U�A�]�Ó��?@^�,D�e��2œ�]	c�1�1O�Sl��)��\ 'ޜ~�|MSJ��Ć[eC�+��� [�H������/$��_�����B��YI��5��o��p�$a�Xh�.0�.A�(��ŤukÚH�E.־_]ڬ��~4�k��
�Ŷ�0N Y�`p�̗������Ӟ��:%�ͫ_���N��"���(�O�>�dA0w���>Z���(�����zY�g6bĎj2|�Y�i%dc���oJ�[c4�N��UW�h���5`A��}�0�&�� \��J C����=,��=nߩ�
�E�=7�t�J'\��:�����fW����k����+�s]L����TR<�J�QB�7�%��`���v㵛�5�˨"W�X�t����B�ncJ7آ��oPu[4N"$|u�>�?�;�.`��`�
���}�X����e�J$��uN�`�z9��Op��lʪ�p���!( �'d`c	��[���ӍN�ǭK�L;�۳]�(��/�)��s�o�&���a_�����)���da�����r���aV�&�����ve�BU�X�.���$�=%�
zn�1?�J��`E(��aRQ��fjmp�	JS9O$Q���E}����N��^�%�����c��IJ#��>	�������y}�6UH۵�y�F�oc�r�"��~D����>�Č�KW7u�G��i2�&�^��t�Nzf&�����aW�[��g#Tݲe��2P�U�6��g5�
zC��5� ��Q�6h��Q�h��}2�9��ߕT"�/u�,�M0������w?fٞ�d�<�q�G��N6�g�U�!_�H�װ=r����sۿ64����h����n�	�]ܻ�:�����ট"��uO
�F�=�3���xE�``�j	+!q��$=�u4����Hv���m�J[([t�p1{^t���#�|=f��e��.Ļ���fe}�HV���x�&쁸N`v��Up%�����_�Ne���a�@W45<Gy
$�,�n�Zu��Dq:.L���0���0u'�������i
���f4�Dm��v ]t	��)�C(�1Jp�=Qg9���g+ր�@ ���p}Ȫ�p+z�2����a�޻����+���s����iEf��3~rHů_*� B��<��v���<b.#٤v1��5��^������]�(2��dW�(�����ҝ�M��IN�0�Z:����r/��]¥ɵ��w��T)A2,��DKB����)���2ɫ�ͯ���:_�|�� g�����Ph�O��G�^b���U��|�Wi_պd7��\���h�B����Q�����MV�T�ƿ!�y����.J�i󖯭������D��Vo����^��*'8��:U�A�	j�;fq�5�PC��LWFo����{&�����iZĹԶ�
���_�^T�Ag���vR���{2^7	XH�/���G����ȵ�å���$oe	���8T����6L0�4�� E��}�8>,tB��|]N��9���#��>;}m�����q�Ӌ��<�Tg�2~1Ĥ�v��q\����Z5�>��p]G������N�i(�{,+1}��-B2{�����1XED�/�lW�~��@n��/��|�1+�ΣQx��*���d.��������"m�j�Z��6�R!�zۜD�:��bH��㥞EqL��l���m~lJ������s�+�p�%�T���bx��Zrć<����)�v���'�JQ{+-���Xb���~����& �L��*fL[q�0�VS�4[m |ڷy�o��i��$9.q�*��Π�f�$�0uST;�G�ҥ�7�XqyEI����/�v*��%��,~�@�a�D�뀢 �$�-Z��(3��3?<�W�A�^R%��d \�&ۙZ����NA�U����(Hv��1}nu�-�b=cfj��G�p$�4y�T�ϴ�v��a��%���3�b`�4�8������K4���|��A����-���~����*�\�绦��'�����O���},�	�������>�Ԛ[u}���F�xF��Ή�tL�1�p���~��{"���QK��"������8�Afy�S}�ԵŁh�A�OO�{4�Vxx�0��	��O$�)Jʊ5Q/��*�&�2������i�NŶ����q<�0j5A%�G*���aUh���;��~��o�S-�"��UY�F
q��e��6.�-���p�C�ޛ��F��6r��{�d܎��qF����5٫}yI�!n�Ԝ�3R
��?���|�y�*ʕ�D�W�G�2Z*�M]�硖y��'��x7��V�UTx&��Hb��	��6�=l�~9J+#y���!5 B.M@�Oz���>�<��"
�z��m#'q���!��y�T4��M��`��kWdGpXfDn��Pѻ���G�İa�
\�A����*�0�]\���R�k��EWΙ�]%_��&�l`�D�������?�K�5(n�Ҷ@u��\@����ޠWQv��c?R�*���a�z�����+5��m؊�|#���\�M��6�}e�,7Ig�j����/`�iK�4,�Ok>Ӓɗ����7�B�����N�E��YY*�
"�80�GB��v^__;
>[G�t�/�W��w�Lcp9����%Ԛ�{���BY��$j�'ۙ.�^E�����+�k�#� �7a�V����v��w�
��49�(��i7q�i�M�W]�
�nޠ�"�6��\{�x%\+C��MQ�����?�G�(���go�Z��i�.������U`&�{,�F����N�fڣLC�d��5�p��sdD�ߝ�%XOL�&;�Q9F���˶9�����bN�C1i�*���+����[qI,��i����!V��ڦSȄZPx|,]{���� 
��6ű?/��a����xk�,�1���r�6ek��cw'��M? /1"d)a�L�X���������!�el�h��QT+/�T'Qdc��D~-a\��S)�Q1(���@X澃O�k_$�G�3�������3� ���D�n����Ɓ�n��;șe��_3��lX���I�&�� ����bC=�2����㔔/EXk��'w\��XŘ�4�<�:�\���MZt��G	iIp��%.�t�)n.7 v9@=D؂l����mBp�U��XD��cG0�<v��Me�L3�;Gi���^,=�H+D�����x�e�s�/��VF���yf~�ifV��^�N��"³�O0�;{����*��2���k]t����^YQ P0L�U��C&�b��b��!��4��м�w����!�p�!k?�lu��l�����0�&�qB�m�y~/b��y^�kn8����L�w�>4�؇R�� `�K{!��e��2�`�R���zk������h���^4�uK9��ô0��4_Ю4i%B�֐KyG�
�����k���^m �UL�B���@x�\��.���f���ܖ5㋣���/;/��-G�>u�)�N=�O�;���"�k76H�`e�#U*�O`"g��=�d��E�P}�Ul=�%��Y
];�﹪��6×�f�?�=]@g����W�q��NxG�D�=u���%�a�qr�g�<sy�6 zj�ִ��r�������GIF�"y&[Q[s��:X�3F� V�u�`$uu]G4*�����E =,.�jK�{vZ��i��Xq�
���S����jg��f���RA�X8������:С���o'J@�@�qo0�u@e��c!k�;&f<�Π�����P���}�K��)F-�����tc�n�'F��j~W�}O�_�����EC-TB]C?����<�Oө�� �Q_�L�{��(�Y�H�;���}*x���e�Da��Q�'<�$�n��?%����v|�࿸\cy� I����Ho9;����3��O�v��#iJ��(m�����H�|R(\~�_F�X��a�����]����b�8��"��r��$�­�W��,�gޣ�����uB��{
�%��hB�s*�����TnG�^�c��_���V��1����	R)���̈́�L��xm�dg��
���fݤ�.���ȍ���n�KU��d[Y���N֓qA/��|��	v~��=@|=��<�"-"��aU9�޵�D�s,�ǽ�A	ѴCN�p�g�u*��M�2ʙ0x�U¢�Q�� q}~���W~��0-�c�Y��1i9F�4�H5�n���f��ߒ,S���,j��
_��r�r���M�3G.��M�7�����&�1���h�cE����\aX��:h�8~�a�q+Ljr���{�E)EQx�*=j���)C�%94cM���c���Hf�Jl�� AN0�C=�s�W�|n Ћ$�����d� 
+��̍��ZɃ����*ra����1�w��G���tl��X�9�c��.X�yٿ�]�\�X��o�j����sJ�Z������`v7�\oF��n�Q�pw�����K���~�8n 
H5��$�)�~���#������[�B�[�<��}0-�l��)���"����s�"��l�<̄��l�<�8���$d�f��Ϛ�3����_�r���U����>a)v�����u���N�$��>~v�<����ٰ�U��
�{�)���v(�?��?�K� ���π�]�����s�l@���O80���Cϲ��Z��Z�l�I;tOku@�8ZV�7c3E���u1�M�Jx5{t��p��t��Z0"�(�s�6SS[M��$td�ϙ���}_%@��J�qv�[%r��ﰼm���=����;T���d]@���׹1D�e~�s��� ��0��Lr$�Qԙ"��ے8�Ly������(�9�J��Y7k�������*@��$dyq��8k_3�;�Je� ������<��h��K���8�tܦ���67�
yIxiU�z5�t)�͔�������:��A�����'H������0(t��LSs	��t��r���������&&�^��G�f������.��f����!��Nm�_�8܎ T�G=�������pe�g���7�J���k�9�'@�*�@�)������e|��r�b�\�L�)�h[�aq��zt^�v���?��:�6S���X�}�mt�DԬ��M��y�TF,;ڠ5cJ�4�$`����k��	
�'r�%����șSa�+�9R�k���״ML��3	�������n.��<t���	,��Ĉ,���Х�9��/;;�K-��8B����L���hw�Ott�����J��U^�gT.���Ep�VU����Fe���jb�8�@�U{��=i�y������S�;_�^$�&�w|�PpjR���
hg����f�nf]��,<yj�}M�Hy��?��W��g�C�g��'W��I#RZx�ƀ��=7N��Ƈ	���J��/���p��
���?�5��E�_*{/Kk�g���;d�#��I~8]������@x�@).U��J{���F��B�Q��Ǖ)�~�E�]W��,c3[]�.8�����*1|`�n���%Lh��׊3OJ@�b��p;��X&n�թ�Ua��1ұ?�,n+�ѕ-��haRR��PN���}�/������J�����5��Gy��(�|E���,���̰p8(��#-(��
S)PX� V�lo�-����)Q�g���'�{!8 �e**K�x�@C��g�g����mALޣ�X��[���8H���nSG5��D?&-C�8�ss�#U�v��Ѳm��c�YF"H�D���m��1��?"��n��#_�6�E;�L��W/���|q��7�K����������,	\&Z��,Ƒ�bm?��,i�n����b����d�.�a:3\���$���Kcߛ�Z@��&��>�c��H^�ʃ�F��]~������^k!����4���lׄ P���C]yT����SEs��5��&ݬ�`6(�(�������Þ���Ȟ �cٵ��#�]ǪQˋ��͓>D�&Q�6��V�v�D���/�+��"	�? f��f����z��<_��^�+ F_gi{���
�^����+�"�N�}_UW���0�/f@}{��F���a��B����v+���+;� �D�5�?�/��ԘDš��݆ i����DKe���� ��4�aŪ�!V�!�\�N^K$
q9zjLY�i5QeBmg®��*��բ����$��t|� L��(B*�Z�_���N��`�������y\G�"7(�8f���<t���_l����#�>~5 ��i�;�zh �F�I/������-���\�����ڠj���Iq�t�,9x;������`�q4e:F����bHG�!zy�D%���++�݂���nA��܏��V���84�V�5a��!��9I^��1��@�)TnC�e3���tހ�����@bXڝ�D�g��=U�VD�D��-��rK�=�>���b�p���*a�ze=���v\����y{������fN�9��=�A��:�[�i�v8�6eô4��Gf�&N5	��U~�T"w�/z���1�D��[ͭɛ%Ct���\=����Wh"�ma}<�A��zC$�NS[k��7����[f�?h�F����"����WY���-K����J&W,u[�d.^&s�i���X|�n7Z1nߘ�pF4G�5=�Nd.0�����'��� |��޶��
�-M8L�#��l��O�iy������*Oy��K���1�3^�s���)�4�r���!A��$�62ӤV���1k����%nv�~6�^�:�f�]���V�:}x���BI�LG���WH��
������&!H�.m&�\g�V�����Y�b�D��A'yi����Ʉ�|!Qf
���.����d�7��k#S0�YjɶCF�13I0K�D��}Q^��Q��L�{=��r��Śbmnb2G�`a��Y� ����\]��s��C�����@?���K��)�Np��%�e��'����z�dW�+Lc=�Q�kh㢨����Cj�<��IN��29�Y��r����םR+�Cj!�b�ZߨI�("ܗ�"O���%��q9���X.��r�H����`à:4���@�C���
B�4�B{���>�BK?@�#�b4��Mt�i�?���E�
2Ny�1��A��0���r{j�'�П�D�{�������M�v��w�6Ȟ�+..>���:��� s:�6>8G��6r��u]�Vg��*}���4)cQ���[(����/�/'��[	��VJd���ֿV����wNh0��D!"F�V�!�ڜ<!���-�f^�vq��P��wή�z�^��ȻIn[n�;��>�<�Q�w��Ո|��J�����MbWhￋ������/�L%����^�!Y��. A���+Ô��pk�k��.�������,\� ��)��`}��n�;����~>�?��P�6�����`�<����wq�������MqW� �~>w�;���-A��|nN�
R"&o¨�� _��FL�Ѡ 
��f`9)�m|G��	n�v>M2Q7:ʅH��Ket_ ���.֮d�dŖ�h"WO\c�~�\��H�j�����:��u�Ȯ�p�,����G�K��:<}
�*�=4���5]��*��Y�����FS�K�K2Z���o���V��>.�9n;tV�3Q���h$`~�Oq���	0�qH�k�G����̰4u��^�I�V���XY�@D��S�MN��q���y��mtc1�`��q_D�/����|'�2�r��,8TJ���V�)���?��V�N�8�����N�@tD�'8�<8qTʞ���9��x}� �a_�n�~��6�s!�j�=6�B,ޥ9�����C�;�	����o������3ޡ�R��%�)�w�ڍ��ip�E�NY__"��54/=�i���,��z�L�@X2�GuEF����J�ѿ�Gos�w�x|hF��d�j7�f/���L���Ju\�� x蒁{����@	b�V�t9�<����Aٔfa��oԇQ�8q�g��]I%��)F�.Ѳ[����7�+�d�Z=�°x=eI���淌tf���rg6��!oV��q#/ǂE���n�nI
n45������H���udY�����2$�v�5Qp��Յ�4���AZ��p�K]��mJYg3EUkݦY^�jµqA��$�b����}��vڟ5���R��+��-�] �h�[��ٟFm�I�#T%���g�aA�|kd��2����Tax��*WZ�,�QA����	>�f�,�֏�-�5e���ϴh��(��=�!ҿ&�R"C���C��u禋Ѳ�'"-��Ġ�9m�����"!Ț�]�]�;��L��;���j����z���,����FX@Me�-�K�~�V0P{�l�4wO�ȥP����G�WL��;NN=��W�"�ƞ"Ҷ�px���]�Q��{������O�+�N�g��ZU7���H^P�R`�V,JC17��<����N� R�|�2���?���L��ԕ�Q���2��u�����Pl[��W�FǱt�|@T��'��3a"�*[�Ż�+���:K㇄Vz2�F�J�2�ZqBG�9>}��@���ș �*�8/��.~��˴�:�{���Woq�Āq�~���,�.Z�g����ag�����l�B����(��cv��u&-��/������Z��<��&�8��l'�$��.���Z.k�[��29i��I;��(zԙ#��(�ſ�%�U��%d��}Y��M�r�D�!�b��1�T�;������O��
���E��94�&AZE��W&���"6�f��T��*�>�:�A��b3�ퟣ�y�gI� �3��/��q����6���?��Nq��8i=#���0.���r����'<c�l��Ǒ��������;��z.I���&=`�-�-��r���i�,���U~�6��cy~q�������b���4���L\��*KN h����yv@��jqW��gA�������(�'�u1�v��ᠵl;�F�	P��+����٧/����՚��Փ����D�p"�`��b��A��?���@��pp7��n(��̓����נ�ϺsT�D����=����!J�$҃��zO�3���+�9~H�o�Z��L����@v�a�l�d������":Z��Ȃ�<���ܦMY,��h<��,Tö��N�fG� ����tuֳ-ǋv͂#e�%<��o�=^�y����v�� eY��˄�(w$�	��K�LE����=t��ULI#��N��=�y��2b�l7��������}��8W"���.�2t�Ǭ��Qqk�q�3�Q��Ic�/�Z����H�<j��Ћ�%��2OUb�rɉ��!�_���2W�(���4�I�i��a���d_����/,v9��<���^P�*�<iӡ0YX3,�E?EAPd���4Swz	g����}p6ˮ����v�=�/�D7�<��I���	H�ɯ�gG�G�m�Xv��H`�+O��qݽ<����%o��_�A�_������6�s���`���"��ݦbq,/\�揤h7�Ml����\A����	��|<��@T�L͵�#���}"��c�1�\rq�Y$ހ�w���	��a]��Ӳ�nE�(�m��ǷLuARR%����_���=�9x8C�q���o@�9�Pk�d4�R��w���O�v_���>�P����4F`��lu�H�z煘p�R�4Q�d2D�(�5���<���ϩk��M���Z���z?�;gk���%�����<9Ȱ�q���4����C�j�o��'�;t����[٨�{�nT*Z�w~5y�k
��=h# n4�&m��}�0�Cg��[w�G)��b�:}���d/Y��U����㭫MF���H͎�e�ӹ5~���_u,����l��ԆϜ=R�/$�,�{^!�@�:S�)~R�����-3C��崒��F�8\~��'�j�=��Vc�a�r TT3cs|S��p�kQJiz�MmX��|F�
]�� ��z��|�����4�GF�� l��bȏU_���!fO��T�T�j�����w/m������i��6ƞ��0�H��ځ����a�:�%��4�+,N��A��
���4�;%�,--�PQ��oo�cv��Ķ��5VHU+`���>]�	=H0�rS+mK��a�C�)�OU���ԑ+��S߭=t�iAsǀ�P����ġ?􎑱�Hcml�N��G�m����K�̄�:�P_�p�#ʚXW���d�{9�n��%d���%|k�p�}c5�	�]��T�˩���g�����d��"���%���v��!�����P�-�p��M
:�.�
�J3�I�|O,y�k��֭��i���h�c��'���������t�;��e陆�5�#��p����{>0����%���0p��&���m��=��dR�̖~��d8{�;ڊ�ŀx3=腞E�E?D<UZ�V�%e�-���[:�)���x~L�$\�6B�K�&|#��Ga2��/65�`�M����d���_�5��"��(��\
��o�9򃔉���ʏ@�%�����F��l@���V���ő�,[��#��r���D;f����ǹ����}B��t�E�AP�z�	��i��'��D�T���#~�\�P�Q�v���6��B	폩Sj^�>�b�-�%^�>A�}�H�ς���<3��(k+���	vIef�`s��H4S�M�ps��TS?�1L��4EY~+'�+����fX�E�����ځ4�����q�Z##��xHT���Or�w%U|CPyJ��&/����+6	���_,\+oct��**{'-ʜ���]=��컉��Kb�o���$��ƃ���
��[D�%Fln)��Cz�4�Yp`�jaM�E�H�������%'�ώF�v�1X.vT�@bG!�k�w����J>𛱯��P��л��G'���������f@�j|Ĉ��e��Q�/�[�V�<悈9�y��*��Ƙ�U�c/|��O�Eյ'u���lFi��s���3�퐫���G@�� Igƛ����ͅ�)Ӏ��P����e�OoGԟ�ytgꍙ�=!�k) X�9Cl�̨@ũմ���d`��)9̓�؉sy�>�n����J��?����b�{%~�j�X��͜1�9�k��ļ.��ž���tP���P��X��oc�B��W�FU��3@؎�h+q�o�hP����?�X8���I3�&�~�O8��`�O�vY_6�p�l��Z|S���κ���g����bm`�b�9�Ο��ßM��6�SU��g��^kW9k9SxV]'x\���'@�@�<T
 �xϪ2�AYu���A��<a�d�>x����Cl8ii|"��J�	Q@k �s�|l����KE���� ��yr�`��Qm(��K��}%�w��e2B�����"��v�Ԏ��I�5���Y�M1B�%|�vr��s��<���I��?�>��Pk����j�t����/��2.�4����Q
�)S�T�KNJL[4G��u�K�t����gq� =%��d�)7��Z(�	B�Gt !�ڊ����x$rHH��J�-�S��ͭ�~W���D[�us���D��2�U9�c1����N<v��z�;�0D*,���X6 81�:�S��u"q~�����2�Zi���49q��(K%v�R�N����s�3,^���28�
ڡU��Li��yײ����W���h@I�4�vU�?��չ��IR$����!^������7������"<M�̢��c߯�ϊs�gc���}�]3��[��v��4��x?���F��&��?YU�G�0�e��k!|i>:�(�˶-��ۦ� g��$��Y��E5��!H�"��]�K�J��Jf'������ѮW'��dT�ܟ\\��<p���(�e��>���{^��o��,K�������,�3;4�頟����{���}Ն��em������ Q�	���B! ]��MX5�����4Ꜵ�Y���S|�#>	�~���p�yk�+5i��%�ݛġْ�a�[���!)�F�	��_�NA�[s��Sc�v����d�GB�T���F�X�F���Q��h��"��ǿh��4���V�3�3|�)~��Z��I�z�xU@��Xs�圶%��;��	���{Z}�M<XP��%#`��sN�L���0�N�c��cFs�� џ��!JGs"l��%����R�����	����M�G��^4�$���ZИ	RD&��Z����N�����$���1`�+��&l��,�v~Р����jc���@��I���D�0a�`@�Zz!k�;�U��ƥ�L\�
��%"�_��p�f�CEM�6y"�������P�3?1�v��]�,��ʘ�d�$�	0�DK����-��N���$��A"Tq\OI=vH�Z5�����'i�{9|�uW/;��k}ytb�.uV�nЌ7�#��gHp��x�<�c�*)����:���Z�&Sf�yW8�9���"h�g����v��wPT����Z��~�t]9��#�0Ϡl�γ5δ�ͫE�ip���,�.�3���!J�����2���.cJL<<]6�_�Qj|���q��_%,�L�bga��`��Ӝ�ճv����bD���:����%�Q��hR!���y�6�]*�3Z��Zt�'����\Lg�Ƥ'�z�����Ff���ér��g�gA����[Uo�(��Q�n��k<��en�Mp��z^=ļ����bS�`F�b���� �j�����:!�z������@+�]�¯C�E|��ik��`Ax����cB�i�Âf���l�n��=�o��R;N���j'����n\��
ub^�X��OF��QUi�$;���A�e�v����E�+?<���3iK�&v
�������ݥ�	�6�Q��
N��A3��o/v��~��j�T����B�/�ˋ�<:fvqw�\2f��U|�Mȟ"�P�A'��������;��K�s�v9`<��j�s�^��An+?'$�K 6:?^�4N�cL#'����Y�B3���&SF��P���[�Dدl쭤������n��20�ͧ>���Vᮅu#����R'�l����Qh��:� ��o��駜�#�ަ�SK���.C����ɍ�GQ�B@��6����2:����
����۪�+�1��4�]�߽�`�gf�=�o���2�4U��0#�a��4Q��>S|��ϟ/S#������|<qq�"�A�O)!�U�q����x���K�JV�~��� �j̅8��B�,{�V��J���Wb�32��3���p1,��,T��p���<��r�_l���8}�����T\��pۗ`p��r��%�0���.G�V��}��zl 4�}����DQ#}O��zd��	P�ʟ�0�)�%(�݄�P�
��l􍊃��t���t��P��=�ɀ�����6Kf2B���3٩��1�I�:���\)\SbK�42P����Y^��k��L:Α�ذ.��?�g|j8*��X����?�x�{������5�W�k)����G����ǥ�h�KR
4}�.���̴�B/��;_��oHI���u��#�$P�1�t�Ȗ�+�������h��.-5�J���ʋ\��þ�^|lY���Q;�΄����%*J%  [� ���8JM�������z��?����[���_o����Nn�*��~��%���Hc殭��2Z�J率��^�e�mv�;>TbA� �N|R�&������CT:��Ŀ
�-��*�8���s�@�4V����M����y��#�n7$�����1����f�����x�v]��b"q�:��<4eQ�ekD{�;���;�ĬaF������%��-�'�B9w�0P<G��3��2W��f�5�5AS�-�
F�~�
�:Nh��#�C��+�.�>��k�C�: \����	��;���A�,���6���	?�p��t��ІP�c����*��`�����6���RahOƧ�<?��KcS�Iol�����H�:e'f�����ݴO��'ZGU�nA���c�B�4���g���I����K:��)�<w�����)��h�[U�ś(�`�}�'rM'��j���2�\~x����N��&��T�ljX�c��8�����߬h��j�/��)�#i/��� ��y��"m�qH�?�	��Jwn�V*@�ר���F�g�o )�g�n�����:�
;�eA�o"�*�]����ӕ��&oE�ZjsΕ��t I��)��j\������3p�4	�Zq���V����ğ*��y�~zIPB6��r�G��li�%���C6«yϘ�ZNfZ���m\��8��iY�r@�T������~��Ձ��s �(��e�������S�y��E�9�E�#�~�㛟��1�)��l�ݨ�sT�{��Ը��V%=�neU���=��&0� k�DA�G��Ȝ�����>��=:Hh����X3�9����hD}�)��U����o���>���G@�6db�i����*n/W꥘%��eϷ�/�J��\�G`�o�y:���^�xG���:!��w�x�d����v*�0'��:v>�K�<;���}�m6��r]����;���i�N�X���kF���!�6	[7�E�؝y�z/�;��C���0���Yn���%8F%���ꥠ��� �~��V�#^�ë�.b���l�`��S41Q�A�!��2Hn�ޢ�;܀G��i>}�QZn�(sՏ�DN�II'��D�N�=xk��)w�?j���ә��`�~��G3�ae��b��F�t���47��R��n�%���bsO-�y��8��]���}mQ�d�6��s�/��b�` x�e�;��b�9�H�wr���^�1B�(�Lزן0s�j�y:e��B��.����J�t����B�������q���C˔�V�ZR�%�h�8} ��$��N�m=�\}�(`�{��#�O���/$N�q���c�H����Q��C�pvb�x)���"�YaUB�m��ٗ�%�C�0����K�0H��hצa_I_ui�1�F�P"{KvR8���mE������\�/>�����F5O��#����fi���n��ed��n�С���ģ���N���'�L6ε\���jmw9y����c��IS&LU2���no�lY�婞�@�1+H�.hC�o��4�~v\5�I,Hr�l\Rv>�!YK�ؗ��Pe$���{�Г;X���y�!��6B�8z��$�Z�Zgg���%0��J�>l�䥂F�����'��2���_v���oz��6�O�9�l>k_
m?�V�/�X�]���"Y�v|����i�-O|R�j^N��m��g��J��B�38�r�@��H#�-��<-� 0�:v��\�w��	�DY�.AE~q��i����n4���p�pI%�q`	����(H3BC�J����I~~�n_� ERe��X�m`��K�!b(&���!h���Ū
����v��cv:�ңi�|�q�Lk`g�{*$T�F�ߜ��,�>�
�f�Ȋ����E��YIzw��aކе9e��&z3�,�,��V%�!^Y�����R�F|��~�������H�rW������ޥ�<Î��ބ�%b7 F��.��ǈF���(4��1��6� -�[۲%]A$!�h-·����.3vӽ��O�����6�TMޔa����{,a��ӕ���^7߹���V��H��)*��rpӚ�&=@o��70�S�,�5I��ly	>����it�a�x@]gw5�r%�������ӝ���A�FC:d�YI冰�M�@��8����j']�<� �2�_���� f,�/�.�ыC��[e��kʲ��
S�����b�f4K}K>
&!v�l���z#pY>�M`�v+�W9S���<w9�G�[`f�-����d�A,�v7�mu��Y<�����j|+4��)4xTg�Y56�u��P:䠥nY�=���6�>������~�����J����֯:�Ӵ~g���o.�#RJ�·�rߒ�I�l ���i��0X&��<a9���,�v
���}'C)ɣCP�/�r�X���]�$ؾ,&���1q�͐��iC�e?횪49���;9�c*n�h��S/x�H�`l�����vy�k�=��u4�� s�
�SP�綡�#�*��]��,eg����b�������?�������7������<�t�Q�>��h�����!7݀���AI_e�'4�͐iN+�nQ�F����f�o8����S����E:�D\�
I'W8�RB�9@��;�WF�@�݁j��%_�q>�yH蟜3\v* ź�����
�O�!�)��.�"���c$���;H��I>�E�O,)�V�c��<f�7j��lɦ�R��2c�V�:��S�#{	�q�ګR�h�>^k�1>�Aɛtk#:]l%t���b��#d"R��A\	��� �9�p"����V ��T	���|OԬ�L����%8ìhsw?�7��J�Cb��D4x��c�Pob��V�D�I��2՛W�uV�z�;��oD�I���B���Z&�p�B�y���5`,�#�t�3�MK�TZ~�Z���NBR$����vjT?�*��S�$�c��	E�*�P�-B�]���9�s�]���?���|�ׇ1?� �]pP�<��@�|r�t���!�)j4GvBk�;�{� ���r�.�=j��ݱ�˩b�H�"�'�7�2�n:�Z�L��J����߼���4��T��Ҝ�Ԫ�u���	�F-bF��1�3!�,����N�~x����L.�zȫ!�>�DB�k�*����ɨ(vu5��n#�X&皌�a�K"X���A�$�b�3�'�L�r}��e�}���o�m�\"&�[8O��d�J^������\��|��y�U�8�,ƃ���_�S8�<'ϰ]�,�Ce�<gԳfזӭ�1�K%���ƙ�}���p���g�e��4�Ñ�j�zA��-��'	C����\V�t$��U��eW�_�q�}v[��6Vm֔��[��iT�[r '�1��
=�w1�!�~4}���)��M���O�X>�*��S�$��M��"��%�|`�b)�խ9��ߍ=�%$iI��riYs `}]f4��6U;���l�̿���dőH��#���̽!�!w�t�p����iRaE��p"k�§�VP�-	�KDM<$����'ʙ!��6��t�l:��T�S���c�Ø�`��t�ø[�2�1L��a��sT�|���퓩[�UȇæӔ7|�$�	��f��_uDUK��n��R�_���T�ȥ_��R��L:%��UN�����MUS��z>�2���y2̫�"3��Գ��đ}Xz�J��wh׭$�&���('`eR�Jx�;�x����W�m�,�MGWD���w%�p~����؍�I}UQ���tb�&�?ݫ����p���Pg��% >?Јa@\�/*�\9���
a�Rj��ƺD� �eI�Vj�q|FkSڃ�rx�n�H���B�'�>�D��)(hf<K�:�^С4g�>�Y�i���m��������:�b�f 5 M~Rn��V������&LVDP��m�1�TeM��6A��׶�NM֏w!�X�{�o��2$�!�io����P˱n�Y�?ِR���E�\��/x�r���:/�x����F�5lMԧ�/Ǣ��?���b�	��/�Aj�t��a��3f�|j�:�
�k� �X����6L�`S�Cf>�Kt+*s��H�Z!�|w�Eq -�9�X�\ld(�p�Þ��Er���v��(�B{���k��MZofEv�@��ogR슸r&��~�W�u�}'Z�/2
��55�Rt'&�j��w3�td��� ".���@�y�n��6�<^<j�J������g2�d����3�K���E�U3�=\����F`��;�.���j@���ʊ3��z{���=�5\���� �/�6����l|�B1�����H�c;ܐ��(�Z���EP�i���H�C�t�h#"�}p�)7E�X=�-�.�Z�����f˶�8�Ē�����B^��~e3 q��+yʲ�����k$��{w��m���℠ �'�O��$�J,"y�B������:2�Mp���I����/��ob
%�]UO�}���M�c�	\��Q�֤.�;H��d?j�5�Y�tm/����
LMD�s�G�J���iA�y*�)�s=&i��c������qT���q�8$B�����I;����Lf��2����eW!��k��~[�"S3�t�|x��g]@'�#��W�Θ�h0��br��X0@�ewԍm���Aע*���2��/�D�Y����$�Z3�-ss/����Y�9J\#%--����-��d'僔�/U%�����Z�w`~�j���%jU�ג�&����E��&���X�a-�M�hJ����e��Jt3b�%>C٫u�4�g�`��ȑ�МJY���z��2cٓF�Y�c����VR4*���퐦|Zꖡ`,-��4�,����c���T�d�9�����V+�H�X)5����VQ�7q����%�� ׈�S?v�)8���X���!�ֻSb�U�
g}�C�Ƃ�Z���C�64����B�W��_8�mu�B��g9���4�9�1�;,q��"a�/Cn81 Η�.պ���]TU��"��_(L#�K�ib{��ruWG�*����r��n��3�ʙ�/��[����\�CK�ȡ-��8����`d��Ԩ�8�X�M��P�X��`���\L����!_=9��1VP\�OR�g�N��Cs:���<0����b�=p]�q�7`����m~�L�v����l����'����~�q$��P����!��a�-s�F̣�J�\�S)-}�2����d�� �D��U3+0}V�ڷ�����ӾC���"jMś��oU���_�Y�"���γ���ă]cj��Y����k-���w�Fq�t�_��ǀӳn���8��-rY�e��Poo�65q>�Ub��\���:X��:�;�bkJ<���[�tky0d���|�8b?P�m��GʭGk��Q̏��o�����C�w[>n��ܛinv;������~�H����_�������'��sU�1�����B�X]u�Uf�S�tI�[6�sZE<�}��$:���TqI�r+�rt�5���đ!Q(�|j��!ӸW6��{�x��Eݛ������ϭ�ʿԷ�'B�������|n^��C��~�${P;ށoى�FA�8��V3ۢL��a;�I�ՠ�7H�k�	@P����?4�Cc6�Q�U$9 ���`����1���C�n�+A7f�cv�r�e�}[�@�x�^Q�E�(�-ǁ[�6�*^ s(�é���Q�e'���ao�tWSk��Oc
~�&�����/'|��"I�>��p���w\G��y��^�5,�{ȷ
����aƑ��o%O}vns^Y��/�I��i��0�v�)7��38r�*vBg(,��T�2-���bS�-�վ7ۑ�5f�{�wv��rojcĦ˗����>m�
�NOZ�D�}�C�ؓ'SU���N�-*/Va�^ ��ƫQ=b���N�rF�����\��"8d�ys*<#�޺I4�9qw�O��J�Q�&n���/慥(����b� M�D5�"�s��RfWʄ^1x��,K`���	}�[}5��YHY3y~��6%��o2�ݽ��ܕ٩�E��+��\�Ę��^��a�Y�Y��9���Y���h�[Z��S�	qi�P��@��c���s`��_\kA�k�U  VB��f����(��lb�ϲ*�a;!��$bC؎J��	Σ��R�ۜ����r�>���&�V�lk��=��hw4�c)G��wٹf�_����t�ggse�3!n�@1�2�,l<�a��Y&��N�5�Cg���M֛4���o�3T���m6�R ݗ��W�7���-����Ӎ��y��CÑ��1f=A������ʽ���P_�2�mEM79F��d:ST^���2�B�C4�{�D@S|PSΡ�Y7�k�BD[k~[n�߭D�h�pX�]M�ܡ��x�:�4�� �xr��x�0�B�^6f�A�v��� !���&���%������B�Fo ($��f^%�>J�q�����M[�a"��fs���+����bR[����N	�g���t?Rr��wm����Pl��uP�)���H��1fL����&�ws����%k?�>_���":-uz�`j��FF.�AZ���h��#��3��B͇�%�>f�`�s���-~�{��$>{G��};v��n��{��@� ���֧�1��;RaNt���T�:��8�ۯ$vy>h�����~��$�j���U��c��桧ٙ�h���z��F�ysG�Ou��uQ}�5���yq{c�ԑ�_��Id�X��;��8��Y3�$��	�HY�K�{��4o}�x`�0ʥ���ӂ�[�_���KW�A�7l2Wp��Ű�9˄o@k*u�1��0�,�Y5��L��oe�q"���{I���#v�<�jXݷ����X"�qB�3�K����	$�"1�4g��e��(���/ݜ�g�̏�q�(kx8[X�5u��n���|��8i�5 �i�����(f��6��J���u���
��w����Y��K➾�Yi�g�P5�1z��0���c:rbn���	���~�U,�-����܌�I��7�?��;�-�*&=2<\j\�]�r6)rO��pN딝����W������o��!�y\a[Mk���M��Ӕ��u`����Vϛۊ#�蓆
�N�[ص?�R^�5BP�����yw1�<z�fŞO�Ǩ33�"z�+`Ժt�24��ѱA}IσF��O��^пe_N�7-l��u����n<^���D�#�r��Nk�\����:����v�qo��)p���%�Pc�-��G����ma��FN��`kă_�z� �~���(�o>/�8[����r�[��N��Te K�P@�H��Z�]%z+�!
F����N\#� ��]*���~�e���tfŵ\�x�ٻ��7y�%'e�ӓW�M�۸r&d�k��|֫�Z0\�0�i���^hԢ��C����1���d�h�C�i�`�/�}U(�Ն7_��y4x��tp�Z�n�B�_�N�a"�[�X)Sy�zG�L7v3Nu�W<���;5�м��W<�S�[��b&+P1Սt�p?�u��&σӝW�V})��~J����]tl\&T>���$؞��Ƹ��2K9��Mtںk6{�+�-~���i��X3�O������
�������3PhZ�XtlS�c]�]�샋LS��^�wn,�:��m�k�"��N�6��>:	��3�������kG<O��A���m-9����RH$#�B!*��F[���$��Md��3}O�����4K��,3�gW��w��]q0.��<5��0���h�-�KC������?��G�ٻ��x!f]��:�}i�k��r��Ew�?��CQ���P�"�Jͣ6�z'�r���;U���le#s�K�bc��?
wc�ҥ�J����?���d݉�ܺ���\��N.�s)O�Ը�Ln�7��4P?�zG~+��f��<��)��;\w���N��`�gk$��_�0�*����.��)�h����~Y��b���QR�|��hZ�Lb�'_�j;�ϲ���&��qh�\`�o�i�1܀�fG���cǁ|�B򉤐�uM?��'.�E �$-�!�kՊm�7���7��v��g�"l?��;����iB�7H��K\��y��A�>�f>��$��_j�����J�v���B�L������n���#�{��w��G(Z�:0F����]l�Q/� ���8��
���^P��שW��Mig@kt-���y�*7���:�O��tF����初7��YRE(y�O�ӵg>|�O�)7��$V}�0�j0c�v!�R�k�le
�n8ޫ�T��q���R�M��w��Գ��T���G�KPt=�����0�=����������yThEX�;�o�:<��\�&��;�`��g'��{s���سd���lR� ��_qbR�.���8�[�~�6����+��s��A�X���?��+h������{�FL����L���������ߕ�}l-WQ�����q����$��~g��nh���k������+T���1i�	J����+A�g�%`��7���]W�:ly��-#9oI� ��(.:.0�~�͟dm*Yߘ�2�m������5����K�*)�n��8%��c��e��u$���"�d�#�"Tl�V���eY�3��#���uA��Sk`ͯc�8���P����8{�k�yA��R ��U`�dL��D����Q %c���Vh�0E�Vq�\v�����(fq���>�T����&g�*n��
��Ɇ�M�u1&!��%�Bx�����Xc}9��S�x#Ώ�e��\��j~6pjU��SD?ڝ�M�˥1�74'���x��$�\?y	.�9�=nw�h3'yE������퓹���3Km�����Q��dt�g>�����~=��c������-�@`؃7FQm(��NJd��<9�[/������4��z_5z��s��zeU.H�U[��ce��2��2m5�*4QG��-�� �����LS�6�)cW�Q+�[z�m�	)/퀂Z�������c�ك�L�oI��7�q��J��l5��i����}�F0{���}Qb�ngWQ��-��O�rc��XCl��)�'C��h��yɌ����s��5о<j����ܢTa��!�EQ��D�ӣ8C"d�^X[�y3K����4��v����+i*pkO�yz8$���%ߝ�;�u!!�ld�y����,�'[��=ifT���>������|�0���t��}�8�2�j�#r�MK�L��`dp֞A�6�&�u�E���x��H�_XBQ���lK��8s�n�!����{�GG�<�Bѹ�#	�IX*
,�o�V�H�= X5ݞ�� {�Q_�ڼ{"������~'<#$i̷�����2s	�[��������7�X�!��.����n67<�<��~�H�%��\�i�PA%,��|�T��y�y�v�
��i9 7y�pd�e�c�Mu��:ġ$��.�$>��,$l�Y�!֠�/�/�l%X�*_��l�ò�A�܄�{����gP,h5�u�'#�����A����7��Ž�32LpH�Tb���_DdS�F�?�"��΁;2�7w�7$B�#E�Thʹ�d��2��0� Z�;�/X�ţF�=*)Ҡ폃0B�l-���(�<��g����D�ʲO:��W��;�@a�ڡ����tܔ�M�[0�b���**l�mr:��(F�B�HH��^��D�j �mᇘ���G����xpu���:ˇ
p����&��gn�c���?g����BEZ욗�T�ȸ�7�i����F���w�de��%�]����ZY���ML�TIb����M�]O��Xs���ӱ���9�=ؿ��L3���)��I�U�}�lZ��Ǒ�9�@�M��%{�i�D���kJ����V�;�kؚ��S4ۊ�e�����8���`��.��wT�)�|�]aʶ!ͻ������bc����!�φ��ʩ6G���������E�����BI���a�e Yd��׉��/�ݧ�׎�0�LAx*���<"��JY"��W��*�_
��)�$�#
�zJ������m ���@<�!کu����U�����1ۣ~�z�;51�)���Ծ��D/�	�9	��;�Zn�ے�c2=�<�o�*Q��W ���X�ڄ_i�m/�yK���\<h��"ԥ��Ť���9|cKs��4�z%�E��!�����+ϋ5�Y�<Y��#mQ��IG�ox< ��ڳ_+i��~#1/��*VR��m���y����&Lb[ۊ��47_ۏ)��-��Ro?iF����W��%�1B��W:vb�d�uҔj�)���*Ge"��"K9dXl���V�?G�7M���8ъ� #}n5�~�C�X:����	#��C��e���0��c蕻�iC�����ci��=����
��Uƚ$��8��?�"�⎴�h 8+齜�W�F(��&_��1�A�bF�7�h�O��� )��Y��;��.hAA����k�[��*/�L��O������Q���5�+������%-%����o_��,�������9������qd�S�)�SZI�A�ۤ:T�Ea�݌f�ǩ|��1�]��u���r��xW��t�>U�	ɹ���3-)97��K�Cz�Bʱ��nM��SU�{=��lP�{縶����-m�^C�����"7{N�r,�Ӈ����6#�Q@�+$1��d ������Ѭ>�y˖[����?5�E��{ͻ�d�޳_Md��lQ��`�
�髎w&.���P�g�g	��
!�Fވ{ftp,ϭM���e���ˁ,N��.5���unp`�/�H�L�u�Omh0��(T.NR��&�k��dw=VaO�����9�/�Ҁ;ΐ� A��td#�u���ԥ.3M�v<	B�t������b��3cW�}~�Ⰲڰ����=tF�i�]>�_h2J�G��`��:�?�����(bNQ�lf���>� �=@� SG�V� ��A�0�q�r1�_W��0��� 4�v�$߆�t���_X�Q�S���ߟ�7* �9kP5��rY�T���~�'V���G��{�q��9�Mo��}�r�|
V�)���aID2������)SGT�6��L���_����-�zN�!YEbd���
cŎ^��^:�g�,�N_	~]�W�e�c,O1�Ԋ�'x�L����7B����	xB.h�]�]���]g\XaP��bnv��cT�rH���v�f�lm�{�m�N�n��4h-�q]uK���`t�C �=�w���>�XD��-�]W�ԋj�䂼��"�R0}�����4�7���~�:���$D�$��-�b����jt�F�LL1g�K��7 ʻ�%��ٶc '�M�RsR0�H�x�Mx^�k��2\�w�&2��w�����W�⃸V�����3��1�)''�ȣh}����hZ 񏂍�/��_���f��?� 2��4�B�`'�)=�=�"����T[����}2{����x����0��V(`�{2,J,����@&��i�oF=����[����g�bٍ���y�������f��r�$��qt'�yd�w*ۂƖ��R
C^��%���
�^-L�B#�Ʊ̪��'b�v�٭�s�.ٹ3<9EZ[ �i$��Z��b�!����9c���+%7.�C��/rb���v_r8�|^u_	��7j�-��kt��C�)�'���V�}��"�>�{�r�w��j/V�%y٤�T`S��=idr'����O��;a2̗���<�M��3{��X�F�bq3�|`Hb��j��$%�LW��;���q O�������A��2�c�z��=y�^{�~�����z��U0�CX�$4��̤8�*G��>�,��'�f�l~Ѥ�FL-F�Ħ����>���ܚ[dtS�M�^%Al�އG�$�}�y��K�R��Q��r�R7�	T}�+;���Tg���)���I`s�J��uj�H����u�4�����C�/.VZT�C#���t�%Vr���+��(��mۆy&�M����{�HGZ�v��ଅ�gdI�����=�Q��[��VU�9H+���3m�7��<w�3�����m��~&?|�4:�s{�����{&���d�Ưѱ,�Jt�u2��/��-î
�\y
C��
E/ok2W\���Vw)5q���0�T�忂�9XL�TCA�P,��~Z\�)z�+� `��%v��\B@���c�Kא:���] �����"VQ>��K��T�NB�\�p$1�M�bS���+W�U���j�ks0�gv�55!��E�J���J����i���Qw�{@��վLq/y��=" ���.����C���� =m��Z7���Y#V��������4�7WAϋ�K�/��W��s4��Ǳɫ>17q���xv�f��NLґu��(��YT@NZ*J�	��|8�@'Z�֡Q��=xt��ThR�~���@��s67�y�t��1���8R���M�Aӥ.�B�L�՘ J8�UT_M+\`/�~oUE)�^.=��]���	��Q@T� Vyl/V9�`����O�quo�)0��Ӡ�a9@�L�I�a��܂�90!���R��=}G��2!q-h��r�ۤ65*Z����k�������c��x���z�0G�M�󵫤p�V,- p�?���jE�9�R �����X؎@�d$=��oH�e\��Tw2��)zp�qC�Ey��R!����K�?=[�aR����G��&�?�f{�W�@��e~r�2�.g�QC�|,g�ԏ�������UM�:4�SpyC�8��;�~��KK��!����V0��P_��D9N����,�GbHP��n��Hm��e���b��Ϗ�]I�<�m�]5��s6��ע��:��t�7��U�"a��1��@���\�ϣU���^�}!�jƁ��8���=�'�1	1���ܱ����Y���8���1����	7���X'�=k�������v��1f1<�x֧�P.X���G�w�p��/ew���2�c�S��va>���`��f$f<��q� ��V�9�k�C�D�P��A�n5�| ���|1Y�9B��F�{�6�%���F�V���1o	��1��پ�#$��W+��X�~�)��N/݋�|�������V1*Y)È���bh��f �a9t}��-�m��Q�=�.�Lk(��-	Aiq��em��Ja&/�8ˀё�7�����:���E$x�|���i��&�:�eo��U}�7�X��'�x��B�W\�.��z�����W������P��9{�=�6d��N�pW<|A���?o4�����pa����Х� ՛;�����5����NUu#��0��6�����&D<�<�m�-�$�/���^y��έ���	��Z_��\&��e&%Pd����/q�ei��]Ok���H��.�����>��J-_r��rk�$����j?LV����݂�
SZ-ls�w,/4�8U�p�� /`���[�'��yi�S�Jj�6t�6; ]=���EE['�Δ�Otܑ�S	�X�p�^����71ȍ����]�_朼d|;��ް]�F>�^��f�Z|�w,��x����o7��?/���l{�{��U�*�L
f�?Y��)����"�ʦ *��CSp%�H��^,f<bf�#\��l��~��&b�+#)l�\������y�6g<��2
��� �|4���R�a)�"	����W�_��)�{�C�Tf���ŧ?�m�oF`�� =�uw�M���K�Nͽ��Z�b1�'u�}t�y����;�@9=�}?;�t�W�(z&��<"�������b���1��"����ۃ=p0c^����e9mDse	#8n>�I�6mCƌ�.�����'�m�.-c�Rqۻ�*ʻ j��(c�v���?p�8;<	�� ڍ����c�qQ������^�g5��|������!v�25�B�5���JU2@��$H��\1/<Z8�ԏ�ݼ岐�U0����+8���N��z�!��O����]n�Z�1m�n����M,`0
�o"4?�W]N�켬��x����zFʆ������+�C�7ZEl���Y��.�~�����j���)]�$�ތ�csov�껄Q��~��o�c��t��סc-�Mb�d���moؕ����jxu���"��<��|ͭ��"�8��uYJ_�WG/�6s�c���Q�4^9���BLLWt����#M�|0i3��g��5�)3
.���h��Р��� ���hΫ�q6~8�b�.oDU;���K�[����X�*^�p�=��7��Fl��e�-�YG��:�,��1!e��D���l�rI��a��tD�ƅ�H�����s'�W�O�ua�f\5᪕�O��W-���(�4�%9.f8�P�}�X��b�@�:|A�BN'���b/�}gE�8-��jj��yQI�ΥU�2�(?b]^L*o}�"�7��kzX����ٶ�
��e��/k	ާU펡]WѦ
[�Ƀa�G5���]�m; ���tpp0A���0�H'��(m�ҕ�4�T#pi1�uF�� �-K&u���0��5�V脼A��C��8�ǳ���t�	˕��W�}�x�:2�O
�C?��F�<#��4 l�(��pF�(4����i�'���8 Dܴ���г�[�*��iܽ����Ԅp�5�Q�S�O٫)(���D(Oաc��\�[���/ �K�����Z� Aj�(M�e�O�KYޗ9�����)te�� �q����R����?+)��/s��$�=Z�.�G�>��	����*)�����_�Y@⿠�qm��$@gl�c]gμy�$X��{�7���Ť�O�Lȣ���`�|�UQ��*�}Ͼ�,�'CV
E��x{ŧ�q�:� l2�����L�)&��=��7��_eV��!,�󎂍# lԦ:�C�OV��F�O\C	R3(_��)h�RC�_�:�@���3�2t�z�i�$<D�y��"�7e&����,�ݝmg����SЩ�/@h�������|�CT)�9�/���]#�ؑ����qY�Ta�Io)ͳ\��d�Rå�~�{�,��P\?�P:���g3�}u�������i���H��r�CKO1`@C�f8Y=&L}���*�i%�U�A�$_k�5B���MM��U/\:᪠�I�^�H0�I�DK�DR���+Kj,�x�L��O�ޏ�B��H�*���#,���z��O�Wz�8w/^I^�ێ�T�����Xs`�I�[P���Y6x�3"�N�KTcM�s�_�l�]�+�f7��mB(]6q��{�	au:��ۜl����b�)G��?̜$��<���FY��/ku���A��V[붢PH���8/N*|v��4��&Y���I.�����*�Գ��*��)=|��S&�{}��e���\���7�G�[HK�pV|������6Y�-5��͖!�'19��#T�^8�Q7)�y�Q�>n�]���`Âc`#����6)�ɩ�l�:@��Ye媚ԭbV�K�W�o�~�^w��3�$3)��*�Yl�)��X�j`P�RĖ%I��\X�kuX�F�!=*����Ӝrȣ�W ]�/kB�8ğM7t4�-�J���U���z Ir*�;�����ҋ��'kz�R����/�yf���扃<=։Ju/�������a&B�az/�zOx�,`B
�0�zv��ѯP�JU�����h�ńB���uu�z��aV��԰-��+������K�>5��nM��z������@a�]��>��3��{v�xR54�9�K6�Jfp�$�m��+J�r�񘪟r�&|�_�õ� �}/�	�j��3��i���h�q�
�b�ō����9��3��X��jh7b�̍�v�Q".������� �1��}JTI��˂�ho�/]����RUa�|�����]�џ+����L���0o����A��3M}AE�K.��R�3A�y���wG���V����v�����Xm�7Hx���A�i�h��C��l���*�Z�%�A;n�p5�<Gz��T~����:
�������z/�х�h��K��������Ç�Ed���mà�ڪ�x�����Ӝ2b�[�����F�����ߊ0S �tٟ#���.�4jCW�#����cS�x�[4h���<���~���ϥ+�\]�6=DqI�S8�|��1�:^&�f�d�-L��q��G��#�ZB	����k��!YVi5"��L���&�<�����`��ǀ�yy�w�����g�b�:כ��Y
"�1Al͈� ��@�hz$�P{NOg�sh�_���ش���`Y|�;#�G�	g��H��Z���N����{�<ۆzs��/#[���n0l_�/��:�?�jd:��0 `�:p���F:��%��������%~i�Q�Ȏ_�*HVۍ��qL�gc�j�JяʢĕVG�m�4,_�&�Yp���՟�kD��s����;ꕛ�J�����ЈG���x��hˀ�����*8�ƀƀ�<��^Aͬ	��+��^]�u!��U��!N�&�M,�n�H9�#vK�TD F��WΦ�Q?h��O�7�"^�0��XrW�"��7�H�����?�)�&�6�ͩ�6��~/�T}����OY���
����ۭ���yd���InnS��j����ч��
"������B�����1����E�L�l����<.T�5���A]*josXUicj�����hIA���G�%_��a4���X�����L�R.��"�6;���H���
����4	ǖ/_�d76�����edֶ/�GSB�zk����t��	+X1�Y����k"s���y ��G*6�vI��e��&�ǔ�uO�������5�@�P��7j��"�3��.i~M���RƇ�䏠F��0��R������� ��Dl�.Bg7������^Nw��lx9�DT�t��c��?�c��5^��4����ǒ�Ѧ-t��s"!��L�Š,���,�������ZjSg2S�Ϧˈ��N��7�#��#��T$2lKY�3������Z��x|$J��Ph]��:]�P]�;���9��1��G�/r�өp"��s��q���&[� �9MIԉ˞%	�8w��ʪ~{�7N�(/?�5¡���3�[��Iq�ϻ�_�+�Q�x%����k�ܐ�S.�S<�jճN>�,-���)g)y@����>#�.?}|�D̀?�s��"I�d��P�l1|w���e��H�������:�!_�'-@U�u�M��>���=�%/��s������e|�W��<5�e�����^Wߴ!ޕ���L%3��\��^��1��(j���kpM]�dq��jH�2�Hv�2-�ڳ�ϰ����V�����HuQ�
T@v��P�Q�����b2h�8�yS�d��.��{ȷ�_T��q@� ?ÄT+ͷ�S�#�]��)MI]�C��h�Z\^�RYڃRU���!��-�Y��pYB6u��k�6�Sd׻0��U���r� s�����p��s�[`�l� �*��y���V\�oC�__�����m�`�hM)�Ч�˱�2��KO��~l%u	ұ�!$,��6��IҊ��Z4/�ã:�8H��v�ל
��� *����^��$��4��2�t�iz~�G���ӹ���ل����߭���3~I�0�n�����M��;�lh\�W=���?��~0R���V)Hy/~>;�������n�:5c�D�O;���e�����������:��a.}ң��ĳ�"d�\P�A��e��+�.��o��F@��cn�V�U��j��� 5q ˀ����Ɗ�\:�2��
<V���g���kJ����q�@r���K�dS��t�d�%k�N�#+���s rI�V/�9B�S,�A��^�&��hVH;�"DXoӦ���	q6?4�ڂ�[���|�D>צ�r�OtDHf�Ds�>T6���j���EB�\���L�o.�xx&��8"��N@&�o����6K���� y��x������"���Ո�AcFV�z���¨4�K-�²��	�W�����}?#��/M���|L���oz�P�0K��P�6���=�M���; ��g��>҂a����ã��nwiS��.Tx����r���&��;�>���l�T�!k��K�w�B�9'�Uz�fr��P=����&`3����%�`�{����s�����_�֍�!�R[@�F�V��f��y
L>��Ǘ?m��������mOQ��A�\�-��ND�Ρ��b���N{HY�����y�}F+k��}v��_C1�|SpI��$��o0�c�3�{�B]���B^�^qM=�ޫw3���>yTv�Ok欷��*W��q��	x}{7#�e�x�(�}΢��M~�Ҥ��$s鞐�rG���^�)@88�<�7�.�RI|E��h��~[G�r�-�D�i�Z�1$�鑰�$���&���e)#[\ ���_h!M�
���b׭A|XȰ]c��Ys�B8�k�g��{&�]��@����.� �^���1sD�>�o�n,��������f4W���?w���3j|~&���_.��|8QDI}�I�5N2V�7����3o� &�	*�6��FiX�ޏK����=�QA�l#����Ó���2{|ey���>��{���t�q7���͎m@Z��f�����]�>J���5�����})�O�Ҕ�e�BMY�tVM�ۊU�Z�{�� ����g[,ҝ=d��r�b�yׂ�����q��\L���Tu��EB[�]�3Q=}�-rB3��x�O�]��R���97�!����;����b~!�$�-��g� Ώ:�»]|,,߇��ݽ򴻚�l��gH���

Jl��(4��8��B��PnEUߗ8�d'�bEB����?6��NN%�<�gW����p4�+�J���R�#��=�c�G='�G.#)�q�)��;�<2g�}�`��Ď!�0�� �]��%�P��l�,�Hl����Л1_�S�0B'�E�Q��/6�����k��=���8 �P���f��
�ؐq�v�޺5b8���Q��ԥt�P0�[βqĵIx!��<�4N�Κi���%NS�i���;#<_4RѢ_�����h����~��]A\ĔV��M�����{�̝�u-|˾��5�� D�Y����|���;{��k >��3Q��V��3�R���@5��uk.�D���'�S��<�f�h��ԏ�H<x1�����s5��K!��㙧�&c`:��%�z��Ȁ���\�;�)�m���p*�;h�S6�����A�Q L-x4ʿj���T9p뚦�M�>/��/؅0�ęG� P2(�̊�A�v�it�d�7q� t`yF1�]p?����(�X
�$ق�-�����歾8!JnY�ʖMs�y: � `��"���c���yO��s�Bƞ�qzH�\d��|�����' >��Dr�=�-U]w��z�n�|p=�"`꿻+[���${�m3Je@`?��������W��h"u<}x�<LX������R~��.���U�ĉ5.�r�o7�ۚ:���۬�ӑs��+�y�!u^#��B�5�b���-��\=ʏE�V�����}>�k0;��3iw��]ͷungF%�Ư	�9��-���|��������*�հG@�?@v6��������ӱ4�G 9�t�8������yM��[xU�a�͙�+?�O�ȖN��N�?0]�
�x��nws�:������Z��*d���s�1��˛y�"�?5��>��y@m��=��@�9��߉��̓_�ߢq���FL3N(�7�"�:���̖K�+Ֆ�r��M�BC����[O��gh"��Ct����p�Q둘��_�3]��$�Q�Қ�����
�x&�@��$tQ���S*��v�d��HJ���r���:�"�D۱����u��J��̷���j! e��%3�AX§��w3����(�*�M���Yx�'X���˅n�Щ�F0/b��,lQ,���������3P�@�����?��x�DQ�h�3��.�����]�o��o?�Oҽ�6��~���Tn�WU>�\��"��
PC�7��e�+�`�y�gT��Df&�`�8��-/^����ޗ����� W�F@�12��H,�]�o�CeC��Oϴ��8��� �֊�3@���v[wŖ,6?�|����\-g^7/�=��fJ7�V�/�k_.nV��ͣt=�#х��������Բ�.4!��X�'�f,�����䭙�2�Em�@G��P�g�[��zB�Q��vÒ��$������IW�W�p�����+G�5��C6x�3�=����UZq�7���q���j�3���������"7�L�+�o����10,ǐ���W��B[qz�34�K������|gc&x�r�m̬�i�V%KɱhW~�6[�U7���i����CS�H�x�9����m�T�Q2�i)
o1�2����qPe^���S^����)�-{p!-�p�K���橺V����/�ƀ�4\!(���=@�A�өum*�83Ud��*��)3�m^����������r��8+؅�����:�c��p5�DRB�T����\t����W�H�QhI- y�J�F��y��=�exHTF��������%ܟh��/�D��[�s4@��}7:;2�7�o���[�]w�I7�����(K��}�����[X�oQ- h	;bPI#��k����H���E� ϭH#3ƭ�~�d~�d�+k��ź|�������6h��2�4M����eR�]�y�"�I-fL1Օ9��ꏱ���1�ϴ1A+W������q�:�	�K\u�o̊��O0?�<�o&�3�U�ѡ�h�%MAe}���b��Vjp��P����A@F�<�QRޠl`�b! Tڱ6v�u=}��L���ñ��1�
�]��s��������V�=�%��"�܏e��ɞ<)�~83�Od�������f�]�n�	ilZ�Ym$MA�Fd(�k�j����~�Ґ��0cM�N?��Y��}	3�sHN�W<[��*A���S�+��G=Ϥ5W�E�d���f"�vS �!-��Ǎ�eoYK����)ra	����6��T(��%YWd+ ���$��z�}i��S��H��� ��(�h��dW�j��2�sΓ�ڂ�8U��'��y nA�j���Ѹe�K��}�Ql�8E��rZ��9���-|M�r��=w=��_a��$��2���d���K�����G��k���+"T��(����Q3�^��ް0���u����f��Ț���CIz�0�q�y�j]�s�Y��r�kX7��0P&w�Y�l�]��+�{��`�C�E�\�����ZvJ-\�]	h	�i��Ox�����`��=!�g�ʈ���O�@�/ �#s�}�O�l�|�(���4���}	\��Y�Dj���qs#��8�p~�F���#���"��[���⨲����Ҷ�t�^�UTdY��O鵈�c�>�m�۝�^)qz��uw�CGD��mj�}���I��)x)����#7A��jB��QAtl���F7!7�zw҄Gͻ!�?{�]x�t�t����e�Bӓ�A63}��F���cu~$��pt�wF�m&�ZG�Dp7�*$�5��WX2��y�~�G�.g
~�� ���րI�rt��]n�`��bq腺����VU���l�R�����4�S'�;����(�Xh����W�z?{����l_�|6�S	�e��L�s��G,{�(�[`/��,�E]1D@��1�+�_�ޕ���Uqɐ����p���4?[��y�5��Q�8���G94���=�*�lz]�F/�jc_��I׈�;]���z��2�\���.��o̟8��u�Gg��Sk� �Yn6����sl��]P��K��J���ǥ��?9��^�q���m��IHj_���oi�]�h[������US趴M�xf�vh"'�Rt!����q�cz�h63CW9F��r�>{������!D�r���.���6Av%��[ɦ�߰�D�T��^��s�Q�4��,O�c��T�]������3t�>m�;BMB��S�As#�����D�ԗVB���I�4\����ilO���B�3��E�����#>��ɥ���
]�<dT�Ɲ�A�aK���Mykl(�8)�P�<gt.�tX���$�x%6l��A�֑Q�_ά�2�w�����_@�x<3�������ĕG�.-�nV�\o{_�9u(���@%8��$�� �H�߶�+-����Hųԏb���_Y��[,5ف�
 �[��ھc�~�LXz?6o;��(���$���C�@��m�#�}���[H�_5��Q0�����ky��.����1�SPlN�������oE��!gƯd���7��ETMۛ���9���?�i�����X`�|��b������	����tT%Y��E�M<ѱl��(ǅ��D��{�z�%���=��T&�_�3�\���u0�ɬs�y�[�la�S�$�m�h
}T8w�`�s�7���-d�',ۂ��ɐ��e�U湯�KO�/y�?���nVKB����V �=+�je�L(y֞��������׵<���R��4��0p7BB�A��C�2Ȯ�Ǡ�ZC%Pj��с��
r�ԗV����y-�#�]�W�: ��4�J��̝i���β������)�t(�4�4熠�l�k�������&��g�+>�z9y8,>.��㽻�Y�;1�bf����]Ƹ�	��cܑ����M�}��׉��T�bH�'���|��bZ���:�����dԊ��Z�GK��jI���R-��员�C��ܵG�:l�������e���/NS�Ĭ	���*a���������n�hRo֩�d�z����+�@��
23����;LRH6l�k���2K�%ؾB��GEj�8��G�E���A}A%��
���(�+?c���.�3�-,F5d�q��#��9#����!�mb��q+�(~^��5�}U�@��t������T��@o����̠�9jҏÈ�1F�@@Q����n7TI4(*���G �A���a�q `B�V ԢQN�O����D��z1�%>���WFE���c!�M�}@)ĨU���mޥG�oйg}o�e �t������ա���+*۞\s���ͻ͂�!��p�K�6�U`P2��BlUr�V�5�oQS�C�v�˷�/B^|���p[�~� H~sB��rr��N�64�zJ!��j�?���8�% �.c:E��*C�-�Ҳ�tk��Ŗ(b��Hʟj�R�*�ԁ����}�r�/?>ڝ�(�$:�����
���Pke��U3N���+jP�גI�GCF#OKP�4I�&2��Pq~�E�Y��aN��P)�.u&�1KU��D�-�����b(� ����x�o��}mw�a$b�n-Lg�Ae��^�pj�z�E�ZF5���&FÝ�G� A�9,ą��|uꍜ� d�g�j����a����Q4ñ�ǆ7 �T#*�{���Co�P��hQ��[Q��8דxC��6<)G��qDh*O�B ��Dq����;K4B�Cw�f�k�Xa��Bc9�ݵ�}	�y����y[
��	�ن�hs���QB�D����B���I@K�/~˴6���2G���Wަs�YF�8��H��^~���h�B+@ˑ�W��)~�h� ����pS�gw҃�����>��˩���M���ɫ�b��_>!UB�KP��+�}��x�.��d�W�5)�B%��ao��6_[j:���(�	���"%&@lzb���|�^��}q~�w�>mS�i�\��c���(� 
�t��P���ơ�5ަ7)�T����"���4�F�M"�����=2�����d��:���A���|��w��N�����G��A7�/oj��XRN�t��\�@�$/�`y"�������{��ϱ->;D>fks@����葍>t}0���<��Ґ��ɔ�X���·�� s��g�7��������h8�\Bw�&�o3��r�d���t���d�dES�躉�q)Z�����邖�E�; �lrو	{�R�����9��'J7�z�6y�?���;T�RPѨf�ܦp�w����΋i���0��@��f~fa4�Z�3���g��T3[�r�d�c�B�[00MϚ�ً|��A�V1��t%bAT��#k�JS�'�Di/CµUܩyS��Ԝ|�8}N��hx� ���$�ɀ�����$��)�Ŀ��X��r�1�%EzY]���h5t��ܲ7?G�DK��)�@�
X�x���1�i,xj.#@�2���|&�.u����6�kh;����_�}��j��4�U�gĸ��>���2�B�U��LC��eQ_e.����X|��ج���{��4]����!�V�H�$���$��E5���M�Bz���s��aĂ!(��?d;�k!���*!�Z&�.{g�ބIws��#<��y�]f�
�M:B�5����78'��i���x���q�5�Eb� s̞;���͆�8&�Tp�W�օI���h�UZ��G�!%�c?c&�bĲ��mXN��Ȓ2�����ކ�mA�f�=5��"�߅i��h�.[�qS�`�ʦ�8=�G��V��6�Io�<�a8��BkF�U�I)�3��Ok�W&L>��(@门��>��cq]%/�]���Y!՗!�}֯K]D�	��ꆈ��l�5l>��]��ew��xߊ�H�_^P!���.+ �^�\b\x@؍2kl���U��������x�� ���^+4!����^�n��[t�����*D"�zh���+�����"U��S"�ĒPpJw�`Ka��֪��~?�tB}�1W��Y�w��CU��pd�t�ra�H��V_t�˜��aVwf76�])�򟁰�u�o\ٞ������*)���qaH�0��j��۵�'�pPp�IU�o��z��\Xzeػ:Ҳ`Y\��%95Y�;����#���:�(�m���6��F�ɍ���ӋA���wP]O�����ǝ1�d�bP�$��nj������=u�]ɋNi��u���_i=i� ���Y��@��o6_ u�J� IP�Ҷ#�c��e=���j^$q�.���x�#���$p��D�ԇ�~����ceHz�݂���DVv��T)���%�wc�CJ�I{�&�d��{���:L@x���������^c'Z���Ja%dbUn��	$�������4ɇ�|�4���'�Mf�2���N.Z���~��Pqն䘊ۼy9�X�9����)�7U�εE�C��#Y)��=��h�L=^�db�c֎�<����#���f�f��YZށ_a$�Fx���/6y>jӄ��Fy�z�%�#e=y\&E>=.	X�P��/6��^�[!����U.a�C�8-�Ō��p��Q���]ŷ������X?5YL��7@�P�V�.9ɒj����?m�
8B��l�h���*��!�
�e���nc����Ȭ��W�Jw�v�«����?һ�BׁU�?a����Q�9����&=�x���E�mғ�%&Ȣ��E�ӕ��uf�.�σ0���2�n���k�(�0���|�!�����FaKvc8xҟ�[SP�-C��?�z��%��|ɨ8z��B4
��"���brV�j�  �Ϛ��^�/�ؕB�-��h�N��7)[��E�5�����AC�MU9��l-��),��0u��#N�(�ƶ�`��z�L��l���7�yúS�х�n�x^�f�cGC��a9�f��-�>�^��l���u�R𗍬.t�bmr�r��r��#]f,b_�"��L��{�M���4R� �Ϊ|=�Д��l�I�Q1G�m�I*�@8�����Q���[ ��_�u��r4������sd��~�T'|�Cc��ө`��3`�;��6����t�_A㼊rH��,��Х�\M ġz����3-�.|�<g�$�J]|����\�j�[$�}���|�o1�y ���d�U� tW���{��F��rޫ�+f4\�i�HP�p13�ib�8�1�G�Q���(���o��_p,W{��Ya�Й�
��6��ܧǄ�0�1ˬ�Q~��X�2����i���C�����
#�*��7�v>?��k��^V�e�i�����I��t������߳�J�g^�S�N��^����`�?mb8��ϼ�@��(���*m���8��j�N{lq{���]����?�i��u9-�\�=��`_s�qZʒ���JJx��~c7��Bа��*�ь#x� ����WiB�~���x���B_~N�)��Vϒq@�+:�1��s�/�E���W����F>J.���?��W �H�x�rڶ��7���w�K)z(�����g��/�X���_kXv�ñ䢝谅V�6��0#�	|����F����izhh8���n�d��kK��o�x/\?��[�Z����?�(<�yn3c��]�I�x�U����׃�ΐ��?�%�WW�aX�G��������@���]��:��բ4BC�3�l̍�g�1�.�١�S��ԁ��C����o��VSvی��E4HAu�������¡�z���"o��6�@����S	�HYD�+H�F�7����z�T�G*}��Vrl������<�w�*�K��b! 
�OB`(u�шwHS{��|Y����>���7S-�"�f�.KF
��L
��j,���A1aoP�T� +�t&�H�'w=�MH�����s[�Zd#:�©�B��NǸ�yM��R����Č�E�5E[G�[�*NP�[E�`z��۸���؜`>z�bR1�ȬPh!�_�������89�֞�D�ʰEM�.%���&cV��8����)�yqj�^T'�i�8�~�~_�DzE����D��8�$��p?���Z�p<�<EH_����o{{���b����(P�+�:��&V��Ub¾���XŬ_�ڃ-��S�Y>g����,��:9�c\���5��dR�}ti���j�7u�
��L�&G
�k��%9�,ޖVņ!4�3��H\U#��O���U}b���Sֽ�ң����m� �s�TBN�<��^��|%<+"g�1�I5B,�/��\���n�숖Lѫ�����Øn��f��gGV�/JFr�cq�s�!��[fҙWQ��?f��b2�N<&��8�vW�?,*|��-��H�t��ő����Ւ#b"�66{�vq�x�b���2��P	<�(�q��\��DV0�v�}] Ie^jz�-΍३%@~y&���%��{����ڳx���p��y<W@��$�B���!ʮI��B2����Pq����u��;{���~�ƫ�H�G�XHqE�3�%	FJy�w�p���xbi2���p��c�O���D�U�x���7V �ؕ2��ė*R�w�|^�g�F+nG{�;���Uj~Y�%����
KAȞ���壡�_xө�����R��y�(�5�+I�w�>tZ*��ƠR���I��!�$�Q�ȷ%��N�����P���Z��J��Td���mk��Soz'R�/-�Xn��%ъ�lzv�8�W�u~�h��+ �c�(3H�����v �C�35��L���[eh[�t������K���p:�sjM�&(I�gy[b�>�FS_����G�e�NN0�|���� v@���3���w���D���2ʊ"�S"2J�V욃�ɿx�ޚ�sp_<�Sg�YMF*�����o��~�2��"Ԭ�$�I�;[E+���gf���Qn�Σm�h��W#.E5��X�&�����Kp�%)=��t�<�	
}���:��]�YU�%�Ʃ:���K^���u���k�y�W������]��֝/?%��@I��hHX�6!&_�)g|ܷg�K$D��p@;�O�=�w�ݾ�)��M�C��Rj�<y̐u)`e�<�5�rJ���H�6�<�~�*:��6V��`N��Y	<bo���Y�i	E�O1M1.(��(�g�j�7�k�t#yN�R�ʐ��b���)q�U�5Dx�bD�/����_�>%��&�?�3=�� �	����4P�F 9`�Ԡ�J��GɍͿ���8�M�QN?9��� d͹$�mǟbC�ݷ%��ZIb�_y|Q/�f�Ɏ�w��T��n�銆��"��bR�ғI�\1No�[e�is��p��J�8�7��7U��錭�	���L#�'*X���4��xY*��<l� ѣW�ɞ�r})4Xk��\w �DKЫm���#c�]=-�@��e=bb�6W�r �>u%���[J�龅>.s���Ͻnŏ~����8� �f�'�j������-B����۵��ϼ�_%�'M�\�8�� _����ٗ�K��2p�Q��O�VO�
;,'�5��녡�]�s�2_��F�� v@Q'ഔ*��A�B��a�Y�g�����JS��_�þU�4g_%��ŝ��fIH�<7���}�/�m�sSi*���P!Şa�f�:�r��2��O����eh
@5�kTo�S�2�a���'�=�Zs%�E��7-�_/O��@ܟ��+�V�D�H��F���m���t������]��kQn�2i�plwܲw�Y>�YȆ�E[�����Ak�_s4�\� B 5����m��o�q�]�-�oQ��/�\�f���x���nca�%��!���{��V��,]��D�a��K���~�u�R�~�b9�'L؃���	��nƧ�;K��X�N&t2g*�yAk��$С+�$�kB�.���5d�ը��y��=C�ɺ)E�f��8^��
��;j���'A�K���=-
���M�Y�����Ԛ0�9|��L�)��F�r|f�C#�~L���!q_�!fM�
�W���/A����8^���q����F�"�[�]�)���H9��B�
+4�Iͭ��Eq@>[�lO���`�
.Jʺ��-kp��|����j�B۟��"62���$��������j^����u�L�~Cv�����Bv�#�X$� �ae�� K�����XWA�FRU1������͈�ec����Tnx��0.K�ǱZ򸩝M�[��S	4Șg�CsgW���b D6� ��f�W�,Q=Ȏ�[��?�5N|[㵜�0�xJ���"Op݋�'6���I�Z_$����o���/�M.��a$)9¢�EY10S��IC�jN��:��#�Y0=��q;4���,���4�Ix�E0�_��$쯖lΜ6��͇a�Y�P?�N������c��ު������@o�[�!w�|>�H���R�'�u<�Z� j��q��0� �����+`��uʫ~���,�5���E�Z���N�����^
�����.��F�,�����5ۺ͕w���Z���K�	�g��?��=o��h1i��q{d�AgJ�(���`��7�����/*�����|f���!d���QK��䲇ۄ��_�ܥ#����Y�h+:	^h��S����5�*='��M��4�A�uL<��)�i6�	s�uT�q.����א�o!�D�1,A���+Vyuh���d�7�r#��DѰ��4�R��S����3��������`�# p�]O��m�K�$4N a�h�h���K����[�2����B��ut=��;5�J��cmi�8�=6��&!����o��ӂ@��4MH�4��q�-Kq�P�T�ڍ�b���<u�O����t�r�y̂�����8���+}[�4,r�i���q@��T�8�C�z��կ���ʪ������m�\�V���1Y/��{��3��i�MZ�6���R_��Wd�%���Wug�Lm��<ܵ������.�>A�0����v,�+��fy�������%�"�zŜ豹-�3� >׸ck,��^�3��mէ3��q�F�n�Ň�]8��vO������6-�\�!.Y&�vK�eu����ד���D&�y(;ؿQ*2?T�F�d���l;�4B���iL& �S4��%Y��O��
S���Dխu�s�=�͖����㰴�Jߩ��\~�<�pAOaG3�K���;�/YDz���,�ƛ8�L D�c��m�P�V!�t}�l�6싒\d�L˳>�,~�H���ޠ�Vw.� �2�x�p_P���S���6a�Ǥ�t��<�~d[>@'0��`������u�Nצ����e]��¡O��>�?��ᝀUB)i�גXЧ��h/+�@lll�������n�OxJҚ�����+�I��!4#:�}�1�5䭌�	@_�*+�y��瘖��9o���OO�4�d����'��./��/ퟝ����/4uu*t�B��A˂.�b`��B?��!���p���J����4�3�Q�;�p/wmd�-�D�Z�/�)�5,�~Ǹ=_�X(�&N�F'��J�蝆`m�m�C\�P۠�"J�������6�?��Uz�#�DѺ�Qu�ڶt��&	��e�?-�df����t7�s\im��(�p�R�FK�e�e��񣞴�� �D��]����9�c������c�o�Ѻ�F�"��v�*ޢ~��Z08�F �pV�r��"~7M�P�-��������sR�QhU�glnE��6�]���ʎ�r����T�o<���Cџ W�W�!a[�3��*�Q ֝���b`�����q�whz곾G'�(�\���4�y|�2|,�0�.i4v~?T��<|H��G?�n����q�}ZOZ�*����@�5;T��?ԋ64%���*Rk�p	�^�t��w���:�cDd��j��(NM)X�L)�q{�2����u�[p�?��`���*¾�B���Q
�Br���@8l��#l�.{>]9���ww���;��Lf����,c(��	�sv���p�F��M�lh�	*��Zƥ�i0���qX�*����ˇ`���8G(�&���{zwy�:��C�>�q���T��?�P�26)O��g�W�8�/�~:��&��7W#:Qδ̿����Bɹ���ц�����R59������ƽ�E����\�=.@��N2���]��V*h:{�@e8K�[�Q/U�)a��t�d�U�J�Q�|�ܱv~��_ӨZ�[`�5Uqv{a�e$�w����S�ߌ�ʲ�/o��_��,Ǚr-�1�'-��cm�,�J���hʉj[�]9<�LMqr����r>Τ5y��Dv( �T�8�@�=�K �σ��X�]�1R������FLn�W@[�W\|>�.6��Ӿ����!lo�`AuEZ�R�P�{`�ozQ���j�뒐��1l��Ƭ�ެ]!������ȃ�@(Bt��c�6m�(�(dߠM���R.��
4NC�O�e�h��w��jGbZ{�I��7-8�c|��W�2�ڱ����x�X�m�s�Wa�= iO�Z�@��b!�:��D+?�.�ΜU�J�jH��6R�37�HY8|q�Z��o�q�q՚�V�f��qr�D����v܄j����l~83A�jS{� ��\�k�¦��R�9ųab�<�C`�M��E���،~~���]���z�RC�[L����X4Y��s��!>r���i#��'�`�� �������;��W!?`�$PR�g���y"B,8����"��!u�oª��Ȗ $Pݯ�f}Y{���?C�Q��~'5oYI�Q7q[��t$V{xZ؁񙂒�>���XX����,�F�:��/\Ap��4{%�Zz$��0FT���I���}����bV%E�>�ఎ��ۂ�i�jJ�Y��&ڽm�o�Mf�lH�g��xO)�c�7��{$>}�޽�ų۬=<���N�����Z�������5�n�> \�Lx�w$}�Y|��x�~�Y@��(���H�A�|D���%�7���P��0��[�׍�O=�'�p(rA�	uLȗ�&��q��0�Ө�3b����	x,1�:���j�s��߻s����^pZ�'ibn|v%8�T��ڸ�nhq�qЕ8���ȅF>�	P�ϣ�u���3���%P�ׄU�?�)���X�1��v�Y���	�C���KE3�F �nn��u�@�M�iP���<�j@�j�L������� j1�Y�ffC+|����<6��{
<ąt�$/�h
��ܰ(/9M�"�lQ+ƊCM<�젠���+� #e�P%N�O�w��А=`c��m���z��"bڋHO�}�ɃN����&��W�(�?�d��ŝ��&M�2���N���Ɍb����?��5�_�����/���h*.�[5�@1-���yػ�vD'��i�|��Sf�Pv2��be�Py�Y�5B�����`e��]@�H�L���?bc�백aT�9P��<A�X�%
ADX�W�_���fI��}gd�[�-GtĠ��m���N�P�����.��ZC����t�śaG����M�vf���}TA̝�,��U�ly�qR�M��T���f���L�ٹ��NJ
�,�P�6�J����}p����
��>(�bCx��*R�L�m�D;��%m���G����֣Z5'����:����X\	[�[���{^�D�d%�w�w�Yp?�n�:�0<�<�@I��V��5E<�¦�������)7<G�P��Y���Aq�l~UxO�+h���V��=�� ��O�ۥ������B�f%F�%<y�%�S�b3����g�k��UJ��a
4n�$��������D$�g�T��?M��*��#�`&1)��r�.8���<�k/���j4��G7:���\���C��.�҃�K>[0\(BֹC��������z�m�J�K�\K?�z_)�B��2ҽ�p��xw�
���GE������վ#�ۧ=;�#s�V����@p���!�t0f����/�)��lh�N�W��9�3F1��F��D�v�+զ�*
x"�������CUQe D�w�m�qdF&��?�ro)��U�b
-���ZϫU�کkr���� ��v=1�c��d�;���l[�n��UڻӃƢ�6�KgVթ�2���cF�6�:'��ˤ���Z��#�C-5�>E�bo��h��Ҳ0{d\.{��Z��\�Y�4نP����f�	�i��t��2X���g���G��3��G�t*�{�V��V�n�l�2Z����ArW-�[_W���\���=_e�B6w5��T�h���n���CZ��>_����:�A�ߪiE	�����O6�?:�Յ�S����� 9$�����	���
t#�6�e�#��C^�rq�f<p4+"�A��)7hc���
�A��ۺ�&��b[VX�3p�X�4����[넆�QuJ�ˑ�]�h2. ��H>9!>�����sz��
�0�뜨�Nu���o��l2p����; GRԸ�+��`W��K4�<�R�k��zWS0&���yDg3Q�~q�|���Ebw���5�@V�8��P�����/�в+ӄ�}��d���+����,�]�������'d�X&'����G$�VE`�!A����]�'NM%_.3#ۘF�x�G�eZf��d(I�R\��e1�,<B�ZO��B?��6�E����
K����������uO���_����2�b�U7���r����L��AŴ�������m)FYp�Z �o,����#�zp!Í�t����6lH�b7�t7B0"1��u5(�t�9�ͅO�q##��y���x;h��D�i��wB�g@�-�Mm�Z�g�;�k)�70�,��Epe��";�yrC:�՛��l{֒����+P�{|�g��@?GCםoE^�N�������p��,�-z:_T�d`A�6��733�l��^px|�e��@�Վ�]��)~<�X�6����+�F$�`�����?D�Z����L÷J�2�0a�r<�y8	i�"敠�Md�;@��S_>,�Ñ���ϸ&���P�m�>1�q��s��q��>���&	_�ap�[�x`_���t�0l^t;�"��й�+����E��	�����Yd��t�¹ᴣ�d��is��!d���w�|t�u��'��2�+����~U�v��9{G�]�1&w\��83����V��)A�9~��@mOSY�w�#<h8��_gi��
����6�vuK��$)�
3��N��D�LŔN]Df�rcN܎�A;��)����ig8���$�.��c�m�M��!��im���l��r,W�M�خ�N ��,�77��V>%'������z �!3���Ѷ�G�����6`p�����f-�rꌏ(U�8��c�Ap�ʄho/����zt���N��LJ\UJ[X%�v��~zCF�9��{�v�g][[�-�~}\�*R��&��4ݜ��ܫy�C�|���eAW�d6}_��`�v_��{g�l����*A�zLh;ƿ����?"c��5��:��5W�D;��3�Y6���?�GgK3Ȓ�q�a����i�l�'���D�a{����a��{�ب1��s���"�s����Lid��:��VAD���	��>07�h���׈��Q��N �[���c��:�tu�a���'��0��D�y@�[��=Z�[�����HU�IN��U��u��{NfI�����M���$�)��7�31'h�+���f�2�ki�����Y>���/��2����6��(�}�Z��WUY|#)9y\8{��Ə4=�09����`B��	��7��1�����#�~mn���W`oR�C��G䶁N���w�nR}/ODI���E�]���:#t����a�v�M�;�ئ���Y>�e�Kt��d���]�R��'؜�$W	5'���4:#��p�a��R?Q�i�5����k��7��:Q�)���oy�$������Mwʬx�[��fQ�(��}h0�_AL���j��Ki�u[�V�*�����U���<�P�왎w��J0Fz�BX m�b�?��ޘ��l�1T\ɛQx�^d2c5�f2��'����̏�V��U�ʱ�cg��	�r1�S"	p��0�v�f�|�u�.>����7�HO�؎�{������f �^�����"T����a�����\�;T��H���
kc�.�91�3�lV��B���4��E���������jm���Ǫ*wd'�1�&����"a��u��y���5͟���I`a$����ܗ�N����L����S�
������qɹ�ެ�>]9��7�ң�F9OI������d�xRӅ�*�9�Ht\]v��GPό��Խ��0�U6��ܨl:�Km�R��C-�# jJ��R#�Qd�?G����(qN���e�t�0
yt�?v|��z;��ʖe���R��A����M�,�m��ʼ�����.���������2��f>��z�WE�,1]$7؁��@��)�/�ڏa_��1�4��\�7Y�m��+���vi�
w��'�ɖ/
J��u��.y[��m ���V���vp0$�fe|���ӗ	G#��h��ފ���V��I'�5�R�(�ϯe��!�6Vӝ��hyW�ػ���c^�Ȉ�ߴ92�w�g�`p��2S�C���*":Icަ+��gB#ߛ�(sh޸`��D��tA�ݹ�ֺ���""*�c+ʥ�&�g���d��tA��������VI1iiр c%������55���U�������+���e*�J��ԙ�p
�i_U�oF���_6Xs�Ζ@��i~e5�<=���G'[\�O��&9�.������ᯁcl��n��5d��l��G�ig�n��6�,�"�̞�"@o�U^�/��1��jK�yB�>M�@�9'�����N4IK�/x�P��MA%>�2,RޚQ�=�EF���
 ��*Xx�>�0̛{�n�Lb�9Z�l��ߪ���x@�>0��-x���ƞ�@����jF#�@�T�u8�$���iN�w[N��u*���K�l����x?w������dq�G�W���!�&tCHg馗�Q���E߁e�c����r�Zf��|2��m�j8��&����Ì����(M�a��&���Wv��b[�#�"���P��;p���T�����P�@�����3����Ԧ�C��é���EB��?T�o\����!����]8RO_�9�
j���m
W3t/�;�I3T��f��X�W��QG���#���<��-]�N���V���kw��2�e��D�f��3sd�w�G���X�;��T��=�[!�ި*P�n�e�Tt T�� �YP���Ր�dڂ�-@+��e� �k���+%%�����J�^9r�� %�ģق�����(�]$�R�ר4s�}��/b�@Ї��,	˄����l�)`���c'gf��7Y�
;H��R{kݸ��2c��c��m���� �٬r ��U6��e�:��7J8"e���0��m��/VQ�_N.Hb����K'�}���ڬs$Lə���r'X��]�g˄�i�B��)y��D���榥	3F��_os�JlK�8���ܤL�+�\	A��(�Q�")�Q�:��&ÓN],Pg���6��v�T6@���Z��o��%V�48�*26Q�Q�L�h��D����G��K�1 ��Z�^d=)!m^<�.}kpܚ?�%��2����>�T��Fm� �L�������f�α���n��~�hL'�C)a�,U�	�lY��̭s���D@
N�k�߿��gt������U��LQ��T&�!���ݥ1�����>Z�N��_��P����4|$�8�'ad���X�<��+�9�1�\}���Q�u�2�ї��%+������q�?�v3
��_���ld{r��?>�%HC�����ܰ�d{��+ �:oB�`��e����p��W�`<�D�Ξ ��I�P��<M6�Q#v�uZ���Se)��oC�0Ia�ck|ځmz5=A�y(���4̖X~�!��yU�yޕ���]靗�X�-�4�^��ס�E'�)�UE3�nr׌}��Ƽ��D�$�I;yչ^�1^��o�U�#�w�qs�f��t���>��t;�i�dfl�eV;I-�m
�9
]y'4&��r;Z:ٷ��"�5�Ķ�q����ޞ�ԫ�Q�o����u�FO��N�Z���1L����ڹr(:Ab�gX���r�Sp�6�J>�O�Stv^g+��S��S�lm��U��Ί07�뚷N:���2XWŐV�vQ O#�sV�ym�����'���!L�m�"U#��=�i��mG�����,�V��.�"���th(sخ�'��_�37�F�]�?��]�$�����v�r{��G���=�_ȵ���z��t��U�D�j�I���ĀB��Mc^�D�s_�s�P~M�^��)C�|��N�3&�`���g��3$)�RN"�|�,�"l|ph���w��c
���̀��&���Ħ��9-�Z�	���!�	ş���x4/\&!�l�Ő�n��)IɗxqFkL�� ~K9,A6��nf�����~H[�X�:b���3F;9qp�TPڨR�}��\�on�Lw�aD�	�L@'�F���]Z��H�p
��<�v�:$�l�ӈ�Q��U�4�����[�����\B6�@����P����/FI�<c��^B�۰$Rͱ�5-�����3M�x��/Q���mD#h� ����ȑ���Z��s�19�����>F �u���=-�i(\�.W͋~�Hn'�N*���Y��f�Y;ޗ }E�o���Ac��Y� �Y�R�x�@�#~�������5�Uն��͆�5$Z<H$[\�p�ئ���y/�14�r+N��}�r�äYU���ѡ��O���ߏ���s�m#��C�PGʝ��{'��(*�2���Ê��(�{�K�B�i�q�}�����u�w4��D��f2&ȂTvxS]$�4*3��_G-�3��3Z���d�I7x���'�Lx9j{sJ]׹ˢz_�R�mX�P����J�1�.}XyK��*B;s�œF�M�m�cF_��,}\,֧��z*��������.�*U�MFj˿���8�gz��	�������o�:.}������n�+����\��>��x׻�oO�L��x�L,�O��p���;%0" Jw @��s�3�c�:��䔗�˳��R��N�[>���/�͒��u�z$�x��Zf�ئ`z��� �p��Fd�%>u�:|.BOE�(ҨN��z|�ky��	��m���lƇn�ܟ!���S�ٹ򃜭ك��j#
�(?�ٞ�|ݘ������|�U5�r��MHqB\�?`1�����Cs{!�v}����~-9Y�����t240��oV��*R���!�EB��G�0�b�8�h	��.�
����%n�T���2a���D+�g6�M3�Y+�x����R\~��0GX3�d��*�vq�~@7�&�;a�?CE����$�U_"W�$�56��{F� ղܳ(I�:\s�hÊ�ɩ�����T�\y�-L���,`��I���-��{��S��^�������9i��Pa�Ԧn��!�L�*r�=Sp�P�Ū����\U���A���u�?�|��^$������A����~M�y�L�u�;�?�u�a��5��}�t�!��(��Y��9��l��?K\L�7l:�k��vG!�y��1�꣠�q��)Nj���XA+���7��.�瓜�L�kl������K)o���Z2	�0�56��}��C��_�ܚI��*��{n#�̈�B��#Uɶ��H���^O\����,0>b���ui��rT���>j�jN9�m�ݏ��҄]8�Ԝ{��\KD*Pՠ��x�{r(%��Y�W��+	I��E���� T&z�HF�  ��"-8�2���F�a�"D@�����גUH5u�)$�U��2F݇Cm�w�P�����+�a�������g}� (��g� /Ӎ4�����>?<����m���>u3���� B���e���4��hLS����3Yi��w��;��`>y��!r7�ոd�Sb���E&z<��g�Cx"������2 �Q�L$�O��`ɐ���mΜ��W���g�w�D��;t�Ӄ֬#GKJA��]�4V�`�\N|y�ϐV�X� ��edZ����;f�h	����!�����eւ[����'S�.�S��I5l����ʣ����V~ޣ��p�	���X��[���	��MFs��ğ&�ԂWK~�?�!��V)so��~�0��\��S�v��qX}�8#K�ᅏ9��q���}o- @�L�����	�� #g����j2��e�'�.�S3��l���_�{�ƲCWڷ�NԼ��#����L�ӿ�ߓ�ˍ!����T�4�ԛ�G#0�@��z�|��{�b�o�!q�%���7[����J�s���1L��=�~�o��9���4�����s�r�Τ I�>���]�2��~[���*pS�P,E�U�=��dι�"Etv�>�fF�߆^���@ U:~o�謤S-!�E�"��:+^���A���-��{�����ӵY�G&c+�=��d�&��DT8\���6�Ł��G ���g�%�/�c��'h`ʡST�N��4_��xѸ��ē
HאSK��8D�S�l+(���r���A`���P9vQ�V�������D� ?��S��$/�p�$�ښ��; �BD=۩�$�
U屑F�s�ۮc~1�#�ZB&E*"]������}/s�nKJ�R�Qc�4CTj5O�N��]�}�}gߋ�� i��DW��%"�V�i`��XƩ �Wa��߱�bޠ����<Phl2�����'���΂3�%��� ��s5���^l����_[��	����B@�"�KQ�e�OHo�B��C���ʸ|�t��a}����6a��sxTL��s�����D�$r~#��Β��.������,o��o�0���*�@})���̿��p��Q_��9Ј'o�S�t�CP�B�"�=�R��4�H�̜m�B�nf�Y�Y���^����D��;���(M�mR��D��oD\Xܱ��5���4}`���ľ��i�^�5���B@NM��=��Ic�>���z<EEg�u!�ݾPH�t���h�b�Xzѽ���
�il�S��>0I��%+G�:⑹˿����Lύ��:ȇ�TR�6��$�g;�y��a�U�!%#�w����>�Ź�'�2�xo�?�~�E*��t�IQ�����*^�vg�Z���Ny��r�љ���urB͜��e�Q��cx8 8@�'���j����/4WV)���ƃ~+�)M�;��{�2����o�����&	jd|S��)Wx��̂��O�R�L���Yr�l��=��g=���C�<!^g J��~rmk��~�#���˅���b�42��	d���VIa��hD�v�@ym2����zܷ�c����ͫ.����P�|M��,�������x,C0	�v�ls֥��4��Q4���T��H7���H���d��oX�J.=��>Ȇ�f���݈;��0v�a�(�l����A��@0�vq����d� ���} ���We����a4X2J�c�Rh��#$�k�p��N��$����]t��	xa�ӟ�JM� :�$�$�ǛE2�Y��`���6���lPDo��L�=��#��{�W���M�8����ޏ��8r�a:0F�l�:�a�yK�UKu�-�w� ��m��Dz�ìp��Y��2@Ӧ��@��?S��`}=yM-�ˁ�`�%H��O�8�������\}�5��ޅ� �VѾ�,f�D��o�3V��O��2=]T��NG�ǡ9��veS�=<S�z�tt�������`�e=G���c��?��F��JᏌa��&��#��kȾ� �ۂM�F���P��6z]+���y�]=O�	���E��pje�ةɑ����a�lI��&WV$rِ��8+�	5��!wV/��		IP�s�u/5�w��C������$�ɠ�ǂ����a1}*�Kq��(u��\�[�"�?
o�������':yJZ�N��^�@FX��P�f�W�¶��VQ0:�Ol2��K7�i�뀀Eߔ��13/��n�hy�3���\;7��>��|��J��g�+ğ��� �W�*�7	�xb��B/�V�l�cX~fC2/$���%F�$��tg
a�,&"Q0,�j,����
p��-�$Bz�f�:褣^MT@;�k�D�Q�	��'�IzA���v���F�54t"�5l��s��Y�������G�l�pv�NG�#���))��K�3�FU}PF��VM
/ᣜzh�JF�pd�t_����{�Y'���ɋ���C��-3Q���C�BA� �%j*�Ş�ҷ{�)C�;�E���^�$b�,� ���(��fZƃA�h!�~�!�"G����߳h.�c�Ug��'L'o�ؠ����k�{#x4��)�^wUs(5�&����HJ�P���&.l�rɔ�
���퓋��B|��;���2e�F���r��*w����w����V�_�IW(�d�O:�Cn���k�	�,<��$G��:�l�d�)��B�yJxX��Lk��>cҦ3J���/���u�QHQ�H�dz�V5cT�)����󒴤���im�3e��r��ok����Uo�
}�Q��2f#@nL)���������7�.&�x��%�!MJ���c�&xxQ���� ����������	r���D�=� GAj!y��9\��5��3��`V�4&��;(�jS�W#����x���LM���3�F���(�Kɽ��5x��c�[�V>�����n�dx �k�8�Ȝ�x���J �������L���"��_�4�V�/��D��P�5O������@�IS��ǀ�.�ѻF���
�
w����@A�{61:_֒Hb��j?������'��m�M��2o�"��W�`�x��N�KB=Բ���� �
8\����ٜ�gӌ`Ѡ�Q�	"��/����AiQJa�:�k�U�[�g�<��Cs2�j�7_���$g.�8�$5���n=Əj+�����lQ���S���3��ߎ��Y���<�>g �|�GS�5�SvZ��V9�o\��=�ZZs��t�ق_Q"�T���� hv����1)UT�;�\6�xS��5,�:QǴN���ݷ�+�)!���5,�â|�"��S�%���QIy>J�0���d����gm��u�M��=S%�`FS�i"x��^�Cu�aA����Ji�wd�u8��^sB�� ��B^�#�)�>$_�E��K�����g�_!a}�A���!D�L�kēxz�*fBg	�Dp�h�D���g'���?�f�v�#3�?A!F�o�r��F���m�H��9�B�8xz���T`a��a�ˇ�V��5^	"7��D$�@{y�.e��P#�&Y��,�|�ERk�/�Ay�6�6�_G(`Ih���`�zhܙ+ ��f|�z���M�Յ��5���J���!#(̹�AK~��ˬ6TQCЫ�z��4	쓑:ڵ�~�;�Fۨ �6�V� ��j��s�%��r�Еtմ7��	�N �r������|�UX���~��7�d;��T(�)���Vbx�^øM�u&�E��L�x�b�����N�����dR37���`)�J4�&�Zc����wQA�MY�oPB^����z7}z�?��C&�`ía��Z[1q�._w�>����0K�0�z����y�
`&xG	����F����_�I�|�*���n-ё<����[~�W^|���CFu���]��G�Y�t�Փ}ܱ��a���M�I}\�a̦��n}�Ix9���t(]��y��t۹����n���I#�!���FF�V����4T`��О��zT����s��u>;Lj%礆fi��>�{���>���]W]�R�/�V��WKB�˶\œ\�"�;�p����f�,h��H�%)��в�Xx�u�j9��Z�dyl︆w�C�E�1g��_�<^l�fޮ�W���b'��d�$��s[�,��}Enl��e�7�X9�և�/t"��[��g�0V>J*�@	�S���r�
��I�����3 ��d�$R���~��/�R��j��ʏ��`����L�+���Z9�VX��}��iO��&U�����3��Y#�/X��^���i����f��3TC @|2��&g�_�y�fMQ�>�������hQ��o'�$й�H�³qD6R�h�\��K���������{�M!�݊=��#��4A���5�1��p�X�.���#�~6.9��?D��&��z�DV��Sq��x�q@N���� =��K�+����T�v\B�Xӹ<--(��Qi���3�iI�z5�= 8�ǡ��Zϝ���b�:o�s���T	��8��]IfM
%�d����r��)�0�	n��9I�,�*�I�!���
�0y����+zlq�p�����
U�3
9k��X��l40�J��N!8�&�b��7W��&���*�Wj��ˎ�+����z���,�#Qh(q>��� B�������ʻ���:9�H��� ���Gu}������s�
�Z��u�"C �`���jt��n��Д<�$.����_kN�t�R�O:�;)d�rr�dL4h37^փ�xrN��6 �It;J�vg�Z.I�^mG34H�.@6�m6��G#��-�)���]uY���M����qM?`߁An���O�i �4�k���|o�o����ؑɼ3A���<Z3�y�r�2�Ġ����('��U���ڋ���K����t���`�Wo���cC�8��2j����%���BK�$"X�@��b��t&��lXz�¢�6����1�>��l������B��>8�c�����w��nQl�{��v�"@�5ǩ��Ar�rUך	�{��|��˻�#�!;���ě�I�C�]����,t�]��r�"�)�����^��M�7��(��c�\�5	<�d���R ��]B�$�����$LA�6�T�a�s@^QQ�̔��#L�E�Zw��Dh�s�Ln�y,�B�/����/t�vT��РADd���� ����hN%��(U��>�4�}�t5bV�����$L-����G1(~׿ �G�~�^�Ng�Js�^"��{oBmBА� D����A�p���bq��U����te�U�b��%ӿ?�Qu�W������xd�D阋!�I���F3����KلQ�̏�����0�yt��(ｾ�_IM�i�_���&_͝�y����/p�W�oa?�̞U.@�7���G�L��nY�4�ҕC@�N��`t�O�Oq���� � RJ �'ߒ�9ӝ�KU���.�q3Ǧއ�ƬR��Z��X5�����`�A�'�l�DLd�8��ng�Lmy}eI5�)}���[���u^�5�d;���Wٹ�7Nm�����I'}�P0�;1?�ڡ��H�4�ﮡ�y�N74
�(�y�m���l<g�05�Vt��|uλgьI���NK���TAv�,m.Æa�z���g����!��T��M��
�!�J�D�]��g�%ۀ�eFHW����4��� #�cO���a��Ѕ��c�_�aזˆo���Wp���ʆ�Ϻ*��׮t������k?	C��	{�h��L���Q⿹R�y��X�'`��zp�b����yCP�ݨ��*UbN�����z���΃^��M����N��Ih�]�:C���u��>4�߈�7��3 <�q�����0|:��P/�x�4�k{hp uW{���oyg1�W�:GGRN������?�hI�����ִ^iS&e1�^�d!�o9@ܬS�YpZ��;V����Ҟ�>��lg�B"�_�3K�s��4�X⏒?�F	R`�DH�v�2������E��8W�Q}�ep�YA�-�4�@w@��f�޸lZ��w66��U9࢈˳=�|�D�?ʆ����f.2j58��2ka�7��h��=f���PP�H�]A�p<"������{�����<fׁ���]��pD���izq���~v��S��i\��oP��E���n�,Wh� +�E��%��}���;#b��!��Z`�a2UX7�Θ�b�,��̂j���#h	wχ���7�Z�C�;��"��0{p� �C��ŋ&$����������!��$�	����J��@�|�o�`�a؜=��9�t��{gn�3��J�k-5�y2����wx�1R�j^P�fm�Tv�mc���p����d��X-��`�����k�dF��P1B$�v'���Mڠ��d���DkY���?���Բ|����1�J��<*V���O��������P���G�?Y{l�{�5{G��6���St�).�7���������O�)��z����'h���+D<h�_#1ޢc@��3\Y0l�̞Oؚ�N��f�c]{ӎ�.>�iK�F�2�}�<��	f�Wk;�M����~�":G��:�h�:=t���f�����P(� �����:�t�e-V@�[�}5t�Pies�
L�R�i�5�y#)G�!�ؙ1X���5�!q^瓪�vi��F��1G/^sZ��
��W��ί��I�H�Y̼�gQF?�v{j��[H�t�;����IաƠ�h�8����fd����"�h�g�;�0)D�L�bE����}s]�WO:�#�VcM���K�b�'ȗ�O}H��!�&Z8���+�F��׀�#�|xz�<�Њ��K*W�|
�*�����Z<��n�n�?Z�S7z��Nd��Ѱv�9���r$[/ֳ�H.��Ｋ�^�MmV,���#�C������У}�Z��֐��]7M�x��c���A�v����E�זŵH� ���&Ez�׏����{��D]���#`Y��,a~��J�V�����<����r�1P{�C=+g�A����MVL�-qP�|WpYu�p+;�2 �w�I'�/���Q�����:�i��c���R���q�P��}���B�꛴�9N�dN,[�͖�Fe�>SQ�Y�
ھ0)(����LQ����՛���Țs
Z�('��s!Ѩ��mspNH���>SR�N$]��r�g;��|Cɩ�b�Ǫ]���=�ex��1q1<6��gFk3kt��o��WQR��?��cGW�#��R�ڨl���2>0´����z�08�#�r�v_C��q����M��J췶Aa�S�`i�u̯$�� ���(�?���<���s�>>�3G񅘴��9�iE�X|��z�dE�D[B�� h��ins�~	����]�^���c���2���Omn��U]8pyru�w��N�{�=>��x�����T���'�E�?T�"v6��ԱsX�e5�$C���E�fd!�����1j�h×�(��e�����ό�i}A�E�_��+����|�mzD�h?o����3g\ ��k����$VG�&F�z���J|��8IOo���Ы1�XM��? �����P���/�����&���䛬s9¢ယ)�q5�yFh��R���&	���zG��F3�	��j��l��z�U�P�-�W\,��o�ޘF��j�H-�m�$��L��b!i�~��?}�2܋wQ���$� k'^Z�χk�hSM�p]�7P���̬"Ti�V=������8�%��������%ꓬ|���H��.DS�+^��t�Y���F�勞�{����
na��\֌�_{?;B�:-��P4@R�ڥ�2j���g3�Өw�5�aJ���m.j�89r�CR���ɼT���x������y��K˪wwX%)��Y��ةr��F��ᤅC1V���Q��k����i�&]��|�_�.q�yZ(�$�ۨ��T��L�{2��>�M��Xn�_:rD���M3��M�BAUv��A���C���E��;�))�b0�NKz�*J�گ�_[Ԛ�oS�Ћӊ��\s��_5��{�5M�0�@x۵������{*���
�6!)=MJvq�p���b���(�.�{�L<7^^-6��,��c8ކ�nq�Te$nRr�ơ���.y?��	*&G�L���&�������ma��C�S��ZwW;����]uU� D{���w;��<��İو9#�vJ�X�����Go��N�2�H����q�{�\J��f f�H�k���i�L=��ܪ\�6���������)9�A�x�-�bU*o�IX)/�*PxK��f�r�q*��?�����	7�����6t�y�]���o��ot�/����ӖS��G�1vH������7/YWm��l�˔%̨��K1ėr+
�^-��%1Ҟ!۟�A{_Y���o�m�s�Ix�$zmf��� ��+B��
e�T��
i�*6����j	�N�Q�f�ֹ9�>wLu�*�����b�D��	�F��I@�����d!~ٺ�k�S0 h��X�7E��Oں�Σ[p@i�g�o4��O�WJ(G{Ү�g� ��e�M�[�����c�ea([�b/>��\�����U�N!th����AF\�z��v� B�D%*����nM�+Vb)Q>�1k��-Ȟ�䓙�Ԟ|J*�YՕ�8��z��a�A`2���PpO���絛G���CB����q�_�X-3�����q�������u���q���1�,�=�d�*�?��m��'��2ɖ#c�L�]���9��*��D��"�j��2��4j@::a����Ab]�U���CX��_"<5�锃��-�_�FUV.���U�`�F� ��D 0�-�].�`�i�t��ߧ�5�5*i3|.0���],xMo�~\<n:�->/��:��a���LN���>e%���Z�+�%x���)�f�&����y4fu�6���	c�7S�C�n�㼅\u���u7�����s-�@��;#��
&C�$����U������˜� U"���4�lci�P��O���pZ�(��q��WLZ�P�UѤ+��̩�ǁԑga��n�L"6)�+��U_���_X����vC(8����D.��铻ӵ��`E��F���>#��2v���؋�i%@�7-f�/^�Hl������'��%�kۭ-0*SF�."o�IE�����Ʋf�H.�j���]�P��?̾�d/G�:9w���;��V�u�@��E�A�>G��ǝ�̐���{k���*�U��
�wA���\�����8��M�t�����A-��o�4Z�k�di�uv���R$�:$yˮ��#<0ּ&�j�H��J�F0-�T3B������O�o��މg�۬�GGq�7��[���7�r�7�^S9={�$���L��#f�:�}S�<����eXW��^LMJ�
V���"��:$/�^�=�����f��~�fs���e����Tq��-3�E�w/�GqUW����-���*{�}.M�ϑ�xA�3��(~ư�q�xp\S�,�Z6���0��,�R����`�L�m�~�ђ�>Wb�Ti�WNZ���=l%J��+h�A��׶{��E���3�z������x�|��+�ٖ���Xd~�ͩI�취
��N������b�F|��m�p�YPMzPG;Іf�ė��@)J�|��|c��V,�b��%P ~<�a:p�X����:�	!b��45����ʵ� �����%|(��ӱ��-·Z��˷��[�`;c�:֋�.=��C|t&+3ʘb�/۸�p��0KPVģ��`�bf	B���\�r�pz�#�8��8����Q�6�c�� ���q,j�������c*�2��Bƥ)��K��9�lHO�3C��%��g�LM���<��:cH|4{��ۣB����K]um��k��J�*b�tW�G�SM��A����>Z"\��2v��Z��K�8���q�;�7����u���O�6F���?�'�K�4ޛ]�xKK��5�Ƒ��������?R����.z��e�\��:��
֗tE���dB�^���J�5��33ϠLB˓r�+��0�M�٫Y�^�i�m'�t�.d�c���3�,Az�l�4��^q#���n`��͇����H~x���A)����}Ҫz�})�o��G��L���Eoy�P�G�4��Rj8������h�r��o�z�>^���J&�@���@Yφ<f/o�t���(�}����5�V�������=MY�be���5('(.*�I��1m���1 I�	�����!O��D���M3k۱�0����D��t�Z��l���>��1Nni57����a����U<N�����nw{bMI�d2u�y�+W���D��
%cM�-�yl�ؠ��	�k�pC�����GV���`�Kg�c#.��|
3�E��KZ�Tځ���m!
ܒo��u��!������k�[��Z�Zj��=�ЋEW'2ͩد�%:��HGu:d�t
�2��4L�����J��^"B`�@�kQk�l1453ѳ�2����[X���c.�I��-3�F���ď��_��5��m%Y�E�ٹ)wb��}@�^�:Ξ.~^���p���e���Y3fg	�w���0�,4М2��W�g�)���g�V8d�H3Q��Ac�I��P����!t�YkrCfJ����V��&�����_�_�J�[
�[+���oHh ��مb���6���aE(H�x��BvҶ�_��'�U�ʀ�8� �u����?����7KF�(7������R�z�q�ڜ��림���T�_��T�֍�R�3>�אbd O�kW�^5�G�-�c�u�(����yzlm8�&�sĳ���.��ڀ���;��@�e�\0�~�*��o��a�<ɑ��䆥�q��?���=U�$!dR��m��S� 񭐎�(�ʗ{��Z��qC�7� ��_��A�&6x��mWt��]��L�����E�\�5���C,�%-EIީ�Ԓ��O�8�#�E��Bə��ޞ�ͷ�lpP4�����^����S�%�  �dRҁ����߃I
��r�3�Tz��%���"�w��᪠XT���L8�PHT�$���Ml�z�M����el2[�K�@�8m�.́
��P��]{H�c�f|�{��"��������|�묻��a�߬_O!Iۥj�(6��}�KI�;��뙥n.�&�+��#A���(��l]\���6SK8��C��d�b����&�h�7�~(|���%V?�mNz��q<P2I�qT��pA-�c�l�H�}�Q��0�p|�����QXŷ��Ȣ�.�f[ԧ�
�7M/��@ ����?z\��a����
,m>�]���������R��߲�Eư���~�'}�������rC��iD��M*sg?��0gp�H�o�@z�[��rÓ��P�U�&��f;�YU����^�OlU4"/��ѿ8��ˣ�8=U:@2�x�a�8&}1!�8���ϧ��!���xCZq8�I����KB�L`C���M�(�-����E&z�+�>O�]U�C�B0IH��I.��\
���c���o=E`�f%J\�_�Ӂu���#r�����Jﱩ�g���>g(�㿴��z_��_oa�>��-���'z�`�!Q'�O�,l!�N@��t���=�D�j �)h��W����u�?�{TLyA?��*נe(�t��M\�Qя�TYO��32�$:�u)��bh����$M�\Uc��,�w��*�e�F0��
P���1��ǀw�L0Z{�(xxK�]mńd��I�߰ef��"6ٳ�tBM��u������\k��}���{��a����{�9��b��r���Lг�sK4Ɠ�-�H�+��#�w�k<���J�P���XgNZ.�q��TR���b �k�`��[�/E�k�G�0i	���@_|�p�=�\tpI�\/�É��5�ؾ��r�hJ�N�V�.�q���2�����iU6'��&ő�5�x�勲QxT���a��M����KH��&!!O�(z�8S�$�C�;s�d�՞UVӌ��i޽���a��[E�e�]�8�W,����e��hd�C�G?�c}FCdX��zX�P����I�2<���kk�zңޜk��-���\$z��{��$���/���	ZdT^˥\�CzL��ۚ V�.�F���hj�6X�a1����G-�V�9�7���'����a�h@�5�g>�����,�<"8�N���P\:cbs0}U�KG�bS�v
�m9�^V��8�B0�=Fh^)���o��וo�f>gD��e��wZ�+�&���ч�؞w��Q(�AP8����p�DP���N��l����k/����U`�i⢍r��9�"�{?*U�:�8F��J(�-x��X��_�Qf� R-��f&.o�)�BԾ�jl=���:)ۤ�/�*���ŕ+#�0�l6�g��؁V�����d��B��E'��+~(�Uϟ�D�����{�Ht�I(��"�v������]0��K� '~e�8
�w�o曫�K6uL2����E]���ؐ=��]zp��WY6o�%Z�`v��۔���ؿ	�c��M~�a��U��/�rew���V>G�=�V���J�4�����UEc�S��c��͛��]e�9,�ru����T2$����}A)0�V���D�ͦ�?�B~�c����B�O�(<3Ks�R������LG�s��=�OA>:4n�E&��B�g�/T��Y-�gK���)6Vi�x>�.a%u40[���V����ʦ�Z���ٜh�Ut�����A�o�'-f.�9��E��Kb�����A7kk�VfI ��O��,~8��_��溺���U�p1�-��0P?:���q g�w�'�X#(��~'ʊ��r�Zs(�P�|;�#�#�;2T��! ڌ��F&�@��D ��C���N���v�TP(?��F���gQG�^��	�-Gy�9��1>Q��80�W�e*k����5�1y#��p ��;�ʶK��JR��}�x\�g����ˑ�td����wE�x;^ŀE��*%�J7W��]��,�rJxIkQ4ҷ4�<��yv����������d��'"ϱ͏$��p�%O����q��E�9��@�hJu:O�v�u����e��v�UH<xF�-����f���%�)��U�B�W��,�M!���ƶ�=Z�.��<������u��|ؠ��!qQր��\��ٖr���]�yj��K�O�lS>����R���w�9(e�:Sڀ��<��8Ϗ1�y�@W)4M@�T `x1Ӆ�bTk�=<�UؚM�T��AMjWrLm�Y����ϧq�)��O�Щ�A&���l�f8gCn���2��#�P初 ވ��B�:�	3i��v(���W�OC��M��3�@�f�K�1ݵ�H����(z�R'h˫�-�靄H���c�m�S9�Vm��L���+���A!<� n$7ѳ,������b�Nq�wM_g���u�����{0�m��Ɉ�z�$NF�/R[	�
��S����u%CP���^=}d�׌A�.+E֨���l�{i�9����Cv����$�G�j��LG�FN�f���Ҙ�crk���iF�s@+��J�-ns5����o��S[:epѐ�"��N�a���&�_l�(YQ?�J�$Њ���Y�O�_����������j��z��s�i,�A	���+��@<�L��o)������1W���-�y�s�����LSy�R$�k)nF�V�P���z�v<bD?���n�Ô1�S��-��@� |]t�B���jOЮ�Y��e �[�I�%�
\}>�H��"���B[���@��H6Ȃ��}x5L%�<j21��\G�K:~����Vq�È���ρ�Eis$��i��nmBtWVƬFaT�４Z�q�¯ҎP�/"�m�̴jS�ů�G���%Z��a��X��qE�9�YȎ��K��ر���*"�1�~��R�2Zs�"^3��j�+��'�L����]�AX5������I�S#k�J����Mx�m�aC�XY�q�n7�N!���?76v�B�9k"&�,O��m5�'��60�r��_Qج��4X���4=��I�f�bW4)�ygbFo�����KB\:���E�3YV�v�ʲN
7��wٽﴰR�W׾��f��	�k�)5t�2����f:@hP�ͳX�9h����aH�<�+v��S�,�{�~�q5�cl�"«H,��X)�p��M�J��U�g
u|i�$i-�^�B�Ot��-�6A�m�A��G��zX���UNC]>�ϐ�.����[ۿ�]©x�6����t���յv�-3�$�5��ҿ)�،t�:Y�(�j7�������w���{��'&=j�?�;����R�|��sLѳn�/T����Q�t�/�����4�F�N��L��4��׶^cӍ˞4؏.I�.�ɝɌ?H�x]g�Uv|�ԄSL��7�>S(ũ�M�+��6L��x�y�����]��=��@�V�'����_ ����P���?�PCҿ��ü��<"�h��%�]�V��G�F�i�̬Bt����r&�x�P ���ݣ*1�]d�ʃ86�"�nA�0V0�,��\q�F@o�*�$ŦĽ�?��F�=?�ݥM��j���w��e��Q	NpZ��B�"�7[q�M��bn+��Y��DI���`�y�Ƨ�k�|��I[[���o����� \2)�&8��ƌ�
�D-	]�?+�' ���ٓ6h�f��] 繯���\�s�1�-P�T� ѱuJ\����>���5�Q~�;�m��:��j�m0�#�=�'l���#>王bJ&'o�3\��?���fP��&X�݃2T�	�v lW*��w�ES8q$W3OA��tZ�|�$Ɖ���vA�DW��O-?��0)2�y4AP��Ĳ���̙�E�O����G�}��+�N�	A� �؎ Tp^�`O�%�����ŏtK�,����jU�d&�)Ӊ���:��47�R�D��X���y:��a]�f�t�SP����i`���m	�qg�c���&S����9�c�T�D�5����B1V�缾οOh�;x'�k`�ώ�/�����Dz��p�w	+�LK����-�Q9�(;�Y�>�����ZXZ��o����`��nP�[�mli��!�y^�V?hN�I ��BV�\m����_���9$5է1}��+Ⴍ�t@�%b�[1���T�67恍s�]*��q��dl�Ř<���N�Hq5�Q&(vx��~�/g/���
�"w��:�7A��J�S�2�����ډ�Ģ&�[$�n�����u�Ho�_�ҕ?H�k���c���#OE"Ÿ`"+�q�$bJj��O�V �^�A2��xd�EUܚN���ƀ��]��<���o[�U�=W�+Z3��c�S%���c;��]�P˵r�	�p��X8���/������z63���J��i�����R�7��\������AI�h`�7ri�:`�
�1��t������X���	Xri�!s��}�.�n������f�4+��Qf݁w*�Hy́�gktq% ��ƀ����q�k��8�����z9�/���k7T]��#��b���!�sm,9��U�����ޭ*0��Ih�oS���*�]�{�=�FO6�Dh������a�Qzvɱ~w�ꜱv_El�GG����H�����I?�ߘB\��iv�%�P��$��v��m�ک,�����,��ýQ�<_��3��+*��@??#�|ò��h���֐���{�����WD��.춉��ߊ�����9P�0��苷+�D�	=N�k�Bm�w�V{�,m�Ơ�(���	���ơa��
+�x`
�Z�Q���Ka��_0�&K����y�" ���
^�@�K|1�1��4�E�[����s*�T����U/l�pw�m|q��1<�c%�7��˘5���2j�b�G�N��Hu�S]�^�~9��f�a�%�������k\����Ax�܄���o�ի�0y!��\t��!��i_y��&�NT�F�uj�K���Z�щ�u:�&�BRw@@�t�"C�Α.���SK|S4���Ch�cJ��?6�q�r5��٘��o)��w?	�� +��M&��]����H�Ĩ1dNIDٙԐ5�a�Yf)'=y�\�qV�`6q �V�[`�CD�fq����P��V�RE�R��������=���,A�9w���֛X!�����١ ��5 ��8����R< �<�Ȗ�1�8��\���Zb_y��S��қ���,�5���x,6��>n���!U��(ԝ�b��|x���=�iZ_l"��<j�$b�1o�.&�ʒ��!ؐ&�Վ�+��:ʦN�7�>LfQ���;��h�*S�J���s/~����ؒ�|M�uD�Ҥ��� ��bMw�8�T	�W#\92���+��+I���H�u�^�?>D_%�zF�_I����l�����&�5��D����B�pe 5E�G�jb���r5��R��^s� P|�� ���\����v�<�t���	2��Wv7K��s
!�l���J�A�?�4���y�}H���9�̝�
#{���/P�Pz6�ЄÒ�m1b*'�tv��:�?����T!�Sl?����o���93��YA5~�v��y
N4'����F~�2��Z�����e���6����L1E4ǐ��Ė�ɴf�r�G)�-[rU��T�~fO�?h��j@Va=�?��Z�u�i�=�|)S�nR4�ZJ�E�k�i�K��ohp;����F1������=	T���(�Cj$@�XI�?$⫗�f
���y2�O��a@��%����]���3'�	��D^�2���J���)i��GNKtlt*��#&��J��CO �v�>��7=к�Y�͖7�-�0�����k��������C?z��M��a<q��M<R�n�J���B;e�e�gV���_Z���F��ӻ�{�$9mF9l��Ӱ�!R���N�(�h��u�"����`��c"��F���0Ƶ:���`&U��3��X�Drob�L����dZ�;k�'>��}��x?���q���p�6 �'k�ȁ-3�RS!��#��(�cS�"�wd��59֛��қ���AiX�;�!��Z�_��C��ӶЂ��tK(����ܑ�ך$��&�/ޫ�VR�E,[���juK(��D��{0BԞ�&Ug"("A?��'C���֛*+u�I����oޡ>�2�%�<a��K�B�|�T��l5�݇�B�X�@% ��9%ս���ӝ`��k�Y�僡d¶�,V�>�69$�9���f������;k�%q�`�����2"����f���}���l�|���R�� ��/�{�!��c�)���.�^q��os��?x��r�JAי}H��i��}>\�(��� >6�|�e+��T�A�Se���w��ӰG���pJ�"-rj����\���E��д��y��02����}7���E�s){�"�)� �V��r�(Ǡ+��l��D�TEr8��tbs���)5̞h%�h0j�a�-�f�}Σ%U����.�da����)�BMF��ن=#��7�v������x�� ��{X�M>$֘D?K<�������+����Ǣy�ҜDX
��k���'��L<�/�p��iuH���������7��}?7R<�J�݄��e�^���',�>���F �D&![�v^�)j:�������jA��p!��;gn��:���j�?J�,!�|���']���� mF6�>H"m/�y:�0����042�a� 93������NWB�[�׸5_#�C�Ї���i���~h���T���R^c��05qm�n�$��`���<��l�����_؂~ro ���w�a2l�_%���|-b��Dd&�T��tW� �̽���=F�R�XA��ڄ{�J3�NA2LU*z� {_��?z�u^F��;5d���ײ�ۏM�����=�zi�;�Ue���~���l>@^h�4��N��bq8�g ��T]���~�{8/e]������0�C%? %�-�����|�5�<�s�*�u� �Vt���Q�=��֏X�/VUT�p=#'�!辠W�Cpm���Tn�?o%�3�$ElJ�l�����4�/���A_���U@��wbL��y�*�����c=�t�T���*�ѣ\f��Ԁ���)DiGjrH�/�@��B��NɗQH�n��5m��fY?8��1���U��8nc�����x7�/U��[ȣ�(A���gL����r^�K�vn8b�Կ6kuR��%-��� a����e+��8����#U�ϋ�#B�����8��۫�@Tc�b�W0_�^��?��!f�1`G�]�%�I,��T���f�i�K��=f�����M�D��l4WՊBldJ� %���0e��W�X��ff��S�Zu�]� {���áC&XT��THB��q��Bf���!��:~��٤�O Gr֝�t�,ϵ�p溑�h�w˯�Wxݝ��ʾJV{�_Ȱw����y�?Tq-������������V�g-@��:��T��x�"j8=�:�E�"�D:u��^�?�0{'���X3\�ۤ(E*/����bDsu��p���|��:���=]gFx����@d�k�}%�.���f�wܾ��i"@wH��Gu���uE
�� ��t=�*������C7؆����p�n��!R���n*u��;h���U ~O\�ڼBR�?==�����?��@�FyzL�9%J>�u��j<%?��[�LhCL�_\���"(�E>�_F!>S�I< ������Tk���'F��N�1Q?Mk"���p���.����>8�u'�N���,E�DM�+�^z�_���u����DӉ�o�	
�m��ՀxZ�����o���vX����|�Ȅ�y�����Gk^�T�"��q��Bp�^tT�����D��緉����}�Q}CG`�wZ;���C9u����5Lq��.�2f~�����M�I�[�EaA�#�LH����Ǿ�-�W��)�h0�U��Dºy�¿0���3dfH��'�O!x��9p��9�t���6��
�V��&�����{��o��PDi��Qe�p���� Nn��G,]ibIߥ"�s��jX�N������z�o|N��+�e#V�	�C�'������� ���xi0�\�ʸ�S}`�H`%��1�h1!tQ\���nb��ʊ�8G�x�kp`ƣ��`q��D��y�|Q��Y�9AgN�b윕@���=��*����ΰڰ�O�	9/�?���0��0���gR��P"�4w�Y!�_nB�S�s\���C48���������������НjZ�r�D)r�^���!�	 ��Z��nPc�,w��s��_͑�&]÷�!}Ra6�LV]�uE��O�"����	"@DM�Ԯ횑Я gj�Ĉ��C����J����&V�"Jv�����ުI�	w�Q�����yp�ٛK&�B2* A����w�"޾�dwuQ�񓣏qb�� 9p� bsv�)>���وݴ��Dsx���<�:�guk�0Wx�[]&�̸�}�Y���	5�"x)򌡛�ٍ2#� ��<׾�H}�஍�����^�\-���p""5e؟7��Knh`��CZ4��iK��7���h�7E�͆S�,���$e�]	����^M+���8����	QU�Z6Y;���ڿv�468�!�O���@��=�o2���,�v��杙����	]�(��^X	�����cﱓW�yo�pK����~H "��΍�}Uǜ'�M3�:	-���ҡrϞHe=Am�wͨ�����ex@1������g�L��Ϫ�O�&*lȶy1�;��Vm��sS�?��6d!�S5f�ٟ:�BgAp�^���{�����������]�� �C˅eSj�"��ryE�1Q۴Vh0A�!w2���i	H[|���)WdO˄�/�vL*�_���Q�lHK?�El͔e����~2��{�!l^u��H���|ښ�":3v-�Ϯ·T��I�)_%��^�l��
��������"H�t�����*�TDc����ۥ��R<(z� ���9R�ӽ�b�[d�,�	GS�79�Y-�d�$+8!���r���tXd��R���b�g�����e5��Yu`��-�LE���5��̣��M;�D�.�W����ޱ+H�����Ђ~����k+�����%�i����B�'5�ץݗ!/��}aM0����0�,�U;�
vո�)[�ڒ^�d�t�㕙�Vi�e���/ӵ��l���ψF���x�5�9j��">�NWe�� ͷR���<��v����"5>�'S���̡�_�q}� Y,�!3qne���ᔖ��*�y�K���F�@�P�x{=o���>��#�6�� �����)+�U��]��`t'�t0�A�����YCG&J���hǱd���H6	q��\��Q=\EQ}�1��?>�deK������H�$MT�[�O9UI���c�&L�{��vBܵ�j~��m~h�+$~c��7@��,�x�2Ԛ5��y��/��y��T?E�׷�G�c��s��G�w���iԚ.������R����Vsk΃B���3��tp(�&���tu�P���/|U��'�@ f�h��(!�b f���g6i{b[�U��g;����7	��#��5��a}K�0H�8A-lq�G��@j����Z�W�K�>KG���o'�{��LaA޿��D4�g��%�0K�o�����W$z�����%2��ao٥O0��T�P=�^����'�	��Y��i��d~?�� �"��{�BuU�

U�=.I�s�Vu?��ZN-Ed�&�e��SA�Qa�(/9uC�(󮃖D���}��6k+	�/�O�}&\���&�� ������$�k���-�Rp�U
^(`4�GزJ�?.~^<&7�e�'�<�����~��\�:0����{iF��
�Ʃ�!O���}��n�|	6%�ܩh`���%qd�n�e�����s#�ž�EEEhΫC��Ó�μ���=e"$&� ͔�ڈM�ºNØCQ����a��-X5�+~D�%"��p3�C�-<�1%�!��9���:L"E��2x��UD��w�����e�m��+(v���/�A�Z�6�k�VVӻy6ˮ* '�u��d�(�E��lWB�<��|�gf.b����Z�8h�?Vm�����l�2�����a �N�ǹ/n_,�r�2VH/��4}cj�aFeEǹ�й)@�|�(��8ʣ���1@�ƈ�$���H��"Oc��m"t��^����9��P)Z1���+�äpkr�	����Q�S�}���&xI[4X[G�KU�埅�3�n�trǒ�`��4�lBb�X�I���͈��|Rf$��T�F|Խ��^)G�����f�*�����A���PDůT�7�t�j��z�	�R.��K����qZ��=���b��4�9*+o,���^u�NX�t�ѩ�Q��5�c_B���7#��!�-$k �5�De)�`���� �*U�@����r��_��eh�C��Y]4=٨2l
�L�� ���	+��c�-�S�4u��>eB횬�ۇ�r�������|t��'��]�"�����m,A�;9]
�\z���d���3��3mL[B2��*���'N�N�(	ۨ���3������,p�L�iA͗.��S�r`]��PLKf/؎��x!C_q#�y�ƜF�!m�7��d�����=�r�y�M��%󠪢V�nɒƘ9��}0�� ����
d�=��7c	
�3+*�{�\��M�\���1ܦu��%Һ��ͫV�i`��%��ˤb3צ���%.%����`��>P��.c�Q9�β��1��M�Vm��H������i�ψ��%~�jy���Buv�O���ļ i�'��H�)6e6A,J	�!F���!郝��&Q��n�΃=^�9�	�O��)�o���5�'Q�Kh�&�@��)S�m�Y\t=���{�B���腳��	��nw���[�J�-� � ̱c&\V���聸˫�۩��T��(�D�5�ӏf������AFm
	(p�c�-*:��y�;ǉ��(�wգ��B�]�W(>R�06�T�9��Gm�b :��0�'1���}#{��e-�?,7xc(�'VU��
�.���֖���&��m���8�]���[y�RR�ѳ]O�x%Y̯1ʰ	��"���{�.K�)�Z�UĢ�B'�*l���5:dv��m@dW�↜K����l��i��d.���)��]�u0z���� gr\�&�r��mD�scy���B�KOu�ap��J桔�Q������œ$B.�x���qz�n���bc0!����?� y�'�+?i|�6(6����tN^�u�*=�S�ع�͇p��e�E}�s<�B���-BM��S8Kn		���e]&��gJ�����͂3 k�bs]�$?���i鉗έ�ţ�K�B�)5Q
'��3]P)�*�Q��4�9����&�P/,�3�˪s�'�%!'8�05�+��C̃���������<#~@�	}T�3�����Ԕrx�EQj���d��1p�b�IaH[:e�W1��w����c9���s��жe��J�q���i��l�<�jo#��^�y�8E[Ɣ+ ^ۯ!����H֓���D����Ws�է�W�,m1�2�b��n��Sz����h�#���W�'7�����E��P0��\\��		�F|d���N��_�kl%e�/"��N.����	zl#���q3�� J�#��O��z�7^O��ׁq���~�K֜#mO�����5Uݰ�zګ'k�f
��g���+��,X�� ��]�gg $���fz,�dgW��n��i��&�z:�u�zF�jЗ��@�:A{:S��0�zS-�F!{�\��yY��� P!�?�>��G^��o-�xJ0.�:�Gv���nR���M�-�B����['d�	Z���>�̿a_ʼK&��*%�:c�,1�;��]��ՠމq��q�md��N����©5cN�/��d����x���e�����^�@_^��w~�ͻ~7��)&��)�m�ڔ��ӿ�ߧ�h��صWv�	�+E[P��7K�HC�]f0)�'g��$�/�Q��$�b�@�]���ỽ�Z���!�O��ٙ_2D6=S��_I?�z�cR>N����͈�T�Z9l��,lϐ��;`�l�|	'��@���u���������R���Q��Iڅ��!Fe@�K�֚�@��i�,֔�p�c0�C��욝$D?c��Q4)u�B�Қ�O�ںQ�W�.�F�����;����C4�] w��[3ra�%k��q�W�_D�Kv�����쎿1-\�e����[t�P����Iy�M-���u��C@_k�2� ��9ǯk��v���d�
��g榕t	�l��٤rL�@�g�-��I7�P�}�^��HTh~}w���*�u<���+�����޴�JG�|[=+���b=uO,g�� ��)C�a����g��}��ު���0��_ I���l�o�2��b�B,�<��J��0�x?-Ļ�N�����Q
�G�U}$�Z�w����i��,z���K`Np^\�_�r���lT�ڌ�A�?�W2�&^,�m��؍ԭc]:�}HbP!�{[l��v9r�e���襌�#�/n�q���i.-�|o �~�3sfc�t�%�Y�>��#�(�{<��{�0���Lh)o��|�Rkg!��x^��VX�
4/��	Hf�ξ)���eمE~紽�$_τ��ߛ��b5�|�_Y�����D\T4;���K݀O�yJZ[���.k$c�=e�)L��pҧ�����|�����iF@���B�2�lBTa#��$q��W�?��(uWV��s��&������7Μ�����(��Qq.�Ash��U�yo�s���V��zQV���ru��=Ce#ϒ��1���TS�X���n��)σ$��@`��W���?,�)ԍ�%K-K��L󭣩WDBe��$�F�+�P0Y&��!4�3:�Y��-4	����'?��r�������ظ���VVjb�Q4н؏�S�$&R�D��G`������ W��"��D �Q�ѷ`6K�d��I�i�FlÐ�����d��r_3D�@�#5����N�����,`�xJ�ĜW����>`[��(&�(��W���t����3eDO=2�<Z�%?�!���	�5rR2�K�-y�Y���;4yi>`,��̧���W����er�E% �\��d,�_,�l�������^��U֏�q^�w�g����B9���O�B?y�I���p>S'#�Cqc=��\�6�J8I#F;.�m�)2Sm�uf���c�U.��k� �|#�R�~6G��u7�q�W�f���ї%P��)��z�AX���Qrx
�U������!n��F�dʙj��!vr�h�v&>��Z��D��B0ӧ�|J1���M�s���Y7��!*ug
7Tl������+F��;��لKz�#��0ni�χ�z*��3�Ǉ���F^3��If8������tffĥwo6�N�p5<�y��xk(н[�?�>eb<?8͌�S"��6��1(l�����9�͊*'���;�k��2JZ�;1�,���s�U�-��P��/ ��}�2���ѹP�)�P���	��rt��Qx�=���nG�~j��;^rw|;���H�Y#��
��Z�>Zѡe��`�O�p����?�!�����Q�ܻ"a�bB��[Ԩ(­��?[H��i̕�T����+�%�5H��c��s���QZ�-�A�G�t2I����1:�vԚ+qE���X�t��H�r����Fv}^�]#�F��������~����L��B���0`�AM�鬗�oA��$ƣ�,���> (ѝ����j>�0�6����}O#b��|ϡ�|�M�S �]��iP��|m�P<�DM�=�BG> �9�p�k�E�܎�I�hC%Xct�7	�C�S7J�w��+Xz7$Ǹ���Iv#�1��{vT��s�yP�4�Y�0��R|�T.�ȣ�ґG�3�����t?9~�_'q^ѾC��y�L�|0VX�A(��8Hy�uR�*W��Ab�/9�v����
ޕ�.�!tT��Y(���9J�;�A�s�����\�E:�#�3p��J��m��F.�.��<�޲�,VD�e����2����$PV߶����Zf������}�4WXV ��)P�
3�O���d0vH./3o>T����ϧ���Yw�����ެ~�Kv�!��Yno����`է2�;di���� ����_	P��n�4/�4D���S$���b��2�Rh��]��a�y!���:�jp��d�4��Ybh�[�k����M?|��XbF��o��v��gJ�X��.ԳC�aD_$��<=���\��r��waN��ĺz)�\%Xݚ�'��:e"����F��#"<�8j�_{�$d���&l֡%U�Bм��)��J��]-vGO�LW����@��}��佞,�a��]B���s�y��h��N]̪O� ��,B���2�!�o?1�= �&PB~�(��l���i!T�U��0f�
Z)R��;Ц��M�i�B��dou�1�wUyo���:�x[n�W�X�4�VF-"`��-�<����Gqy���I���Y�>�;ʜC���~g�l{Lh�P.�Љ�fV�1�j_�I�b�1nܕP&��h5JȊ5�V�z���p�`�D��̬��ۧ�^!2���*[�f3��w�h4�LG֔N#���=�hsJ���Mks��֭/J��7����E��ZX���0�!}���khmކ����.����Qs�w�o�K�D���R;iGx�z����y����9A.���pcl2�ޖ���z�?T����Ջ5�VI�P&�Ĉ��_�
|(<���%���:)�pf�m
�a���%
﫹��i��L��`Q ���}%IT�5 2�>fmk\1:Ӝ���M�3n9�?�ȿ������A*�|��hk���V	J�T->�����O��*��g~�h�3W�
mW C��s�����"a�Q�o+��8ʻ�Vi���V�ρJC������a�M���)�?��C�ߐ�X��d�]=���J￁��j_���ϩ]z��2�
��]@�0�d�߂�-@�(!V�,�F�f�)}�L^[x7�
Q?
c{�#�1��6����|��/#�!�݁_á����-)��n����hԹ�v[���' ��5Ո�� ���w�pa,$N��{Ѱ��-9�+��H8g\F��_���,�B�1}QXC���6]�I<���bkk܇���SI�4�A����Ș�\������/�9��9�i�f�.	�O�<peWH�H�	�fŵrC_��+��%�(���2��	�QA~������:-�Cr��Ѷ����Eys�6��g=�ȡo2�����_H�W�Fx�@g#���F[���ȩ�w�GK���XE՞���y�M��qM �	�\�Sb��������6j.z�y?]b��'!�< <���ǝ�H��1θ�>՜�j��1�0�e��~��Ie:���ruZ�������}�<`X'&��N_ܩ�dp�$|+m�̚Ѐ���l	%��*��C�D%9�Q��[#Fc|��Q�	�W7�I�|�F�_l+�����hc�����^��������(�G�U���e"ju���}���%ܙq�h��s����������|������=�{]A��avt���ٜ}�0�ݧ� &�!pu��)�۹`�2��gH��}�1ި? �ɪ�V`��4C����ӕ��j�TX���2���ʿ�􇿔���ԟ�B=IS1��}TJ&β������]�'E�QZ�v�5�T�7��LXJqţ�ۄ�x�(˺����L�<�"ܓ�^���T!��)A8�ě�_�I�UEY	֔�Op�����~����)�o,}���VU��_ǋTH5�V���	��Rl�V��Ao�������^���=w�s?b<:r�[�B,�Fű�l�������!&;uh��5�&l��1�9}k^��<>_92��a�,�����N�ID�g���$k������Xz�� ��^$�`����nwS	�����~�L�S���&-p��N�<�?RKc�o�h?%p�<�Ά�+���s���&�Mp�NH���K�鬹G�J�� ��8hf$x��(9�A��7��;���������������Βdq�܏��OnȈ$�q�#�l�a#���\e������-x'�R�L�e"�+���(��U��z�Gz�a���s���Ob���5��:!�,d5C^x��x��ۀ�b��L�����d���t�0����cp���r6 `&���?zd���i�2-�L~�43�9�r�=L.��kE�Ӑ�w�-�����qͬ��=k�f�D��Sf�Plx��]����+�p��J��@t����K�,��E�����YR$� �����/_�}��z��A��	�^ �����h�T�=�J�5��n�~��;���E���"]��ÉR��}�nVh���m��$6.H[N�C���L�-�=,S��b�۬{>5-0�%a�|��kfx�L*�k�9ِ�81�vP����PD�@���a�e�Ȉ1*XRo-6��������`�Tr��=��&�X�V��a#{2v������A��e�R��hz*;-/�-B���y�s\��z8��*�[ˆ�	�<m�s�=Hf�Ĩ�;����KH��c��rCR���Ő��v��lDe�ޠW���y.y*O}B�h�� Z�I~��r2뱿a"k=	�=^�{��-�5` ����9�59`�Ğ�vf�I���ug�M�7}��[�	�Jڅ���7G���?<�����qo��z��R���]N� d�d��R��Rh���9�n(��Q��F(������u����*\������o��%&���|	o~�?��26
[�ǳ(+6��ʦCW4+�=Q>�2ꬪ��j1��߲��u��~;Ż�P
=Zv���9>pM�Vzg���2��-�y����4�h-u�aTey	�`��[^��螷�@q�qǌZ+[hX�={�[�L�Ͳ4��S�`�aGX3_3�B��k	H�qE(Z��ޜM%�5�f��<��ƅ���qo��q-�f1��F�'!�4N�*�h�}�5�,<r���H��0�JC�vۃH���ġ��Ϥ�3����\��Z^��im��XS�"�ؽ�Z������B}�����(� d�XY8�%�st_'߲������������lK�k5ӵ7�94VVW�VX]��2�#��/��$h�;��K��AZp@�P0���2���M�&t��"=��So��z���n̲�o�p}�]�9^o���F-�Q
�l��?|kz.���73�[%�á��g�A���7���F��u!"�!�0�lg�*���A��~���A�/��U��nY��M�YGR#��?8�^TE��8�@76��n:�S���R�1/*�+��۷�-,���|]��\�ע!�[�o8��=�����_g�2��U=�f�(t��:�73rD�_�V�/���H��Y�5�{��o�����ux�N��˳��u��%�h�(��}�z������j��Hpԙ���t!;� s$��&&#;#��3�����
�g\Z贉i�u%O����ӧrf@V����w��q�<�_�Jg/��^7+���{s����V�,��r�	���ktgl�z_hR�|@�Skx,_�N˲�ZxYz=�2L���1�X���?��~��r~!d�l^�؋.��ZXL�{��B�a��H��4�k��K�sW}�/4�,|r7ќh�chqk�1��� ft�ω�E
O�
s�!z�'�PW��A���DNZ
�����X��L߉8�*Ж7*$w[v2�{cM,:_֯hU��~��I��$G�?Q���}�IBN�;S`A���7R���d���1U�)��lg���[R��`� G����S�3��>�r����x�$�+������.xB�B;�ݻ��L��Ǜ�"g	]��S����ְ�O�j�C�W�
���':Fds���">U�l�ZQ�n+�9�H4�ұ1�J�����+�����Cs����g���')@#�<��~� K��Wn�9������؏�?���4����+�&C&�t�f��x%q	�Z)߃U��E����Y�x���4{J"�k鳪�'��j�)h+�`�jK�d����3���L���Ĳ韺��2���*�D�^���$r �>��]$S���S�&E;��׃�P�r�"J�L��������09��
�����D��_�O10��he����a�ut�p9�m5��n�$�!a����e�:�8��"�SpN�4 %`�%�7�}��0Q�8��Eu�S1�+�K���x����xۘ��>��@=@�"��� �5�fd�	�Y�Kdz�py��5�|���P��Z���8� ϯa<���c��T;������'tH�����hVɇC��2�d��.� d�e������nWB�L��J��@%m�ͪ�\��:��fo`�w���З�kÉ�x����V|C�ǘ����͖r\{y�g|z2�-��� x��n�4���^����P�į������2R��G�g]̸��u���=z# �r�����Y�O�N�r���"P��:Ş T��R���u����hJ�ȍ+d�?����̊+����EzK��f�9{ cTl*�>Ԩ����V��S��E"�kZ����v�l�Bvz�t��	KE���}�� e�Km�k���R X������{�ć :t�9xFE�~S�}'�rU��P~�|���`5���-�� [}F���B@���$���H�&�hH�;�(-6qL�Z� ]sbx�U���t��v�f<EH��g�``ʪ�I�fS�2,�k�@Syx��-
,C��V�%���9������c���J��OЙ=m�n�@wQ�N4j��?��:K�.2��i��nD��l(��w�u���S'�o3��"�Ex~.�|��m�C�ޓl&[�M���[|� �<� ϵ^ϊ�[�;���w��<�pQx-��U�>��Á�W�U���L��M�40�5eD�����Cl\��!}��N�Y��|T2;���A嶐JuO�*%�UI��'ԒWx9��Cn~��� ����!�ڕ��9�d�A2�Ap �G�,�88�n�R#Z`�Y����")��pI� $�ﵔ0hDQYF��-��
�9����XêT�:��{��{�q_*4�2�(�Jϴ�ف��b#[ݲ�|R���7�Oj��׏�Z���i�UV�����f�'nѳ�DՉ
qF5��~��Ej,6�yf�ՓZ�B�$����8���I�4�W����LjcQ0��Vb���w��yz*�a�An`�f B$5�6���Z����~B���9�Dۡ)�کµ�>�Q��rU��՟¤ ��9�xh�գ�r����v�ޒ6���$�Gu���[��
�;���s�����H��[G ��8��f���a�}����Z����Գ'.`&4n�u,�\�V)���v#�������釋�s T�˻SD�q���?X�r�ӑ�/Y��Kh��_��ҕ�x|�������4�G������N��=��^)�O�ݮ�bA]��z�&,��65̇m�CR2�ј}������j8��o{?ȥ�R������q^������~tԔo�2\�v{޲ �;�
��u�����e�E��R�JQ����g��M]�FY�}Z#@��N<:�� �/�R໠O�'�(���]Z^Wd4��<wq�R#����q��`s��A2,*?]0�w�y�30���9;(&UVkS�:8��v��T-�����.��	gU��W�r���ƞ2��Y�����,����'U�a}�u*������~�ZqiTy�D4��1����x���"�t��׼�H�y&�<BۘU[��!l���	��rݥ����@��y:j,(Lŷ�g��s��H͇�g���=Ϗ��ۀ��2�|(��N�A����&�ُ{H�SÂ|7��f\~$�A�"�"^��
\�[!~HBϓiB:���[^�m2�UOf��*�ȭ@×��A�i�W-j~�N��PL��	!���ot�Qê�8��ڞ��5>�"�qJ�7�4C�s,�F�hc����G�5"�n�n��g�I��z�Q�H�ފ��tH��1��яi��Y��'WS���1���ܡ�E� �󣜸���qI�9-���X8�E?���9��,̰e��+��s�;�K�˅U�i��2���j�����ц}�ֵ���j�~��~� ��Z��w������*10��V)��Hڈ�C{����t�>���*h�E�Ρ$>�ԳR�[�m�v�$�Gz�wRJ�p���+�z��J��
95 �r����ؕw;����&)���_�u�Z궗F�|�1S�\�]���ǟ��z9OD���C��Tdxm/���0�>�P�c��UF�������KYUh�ζ;Ɇ�K�']Ƀ{]d����`w���R�c�w}�i[Q$�����9�����������{Y��W�衁>!�MNr����M"�%�h��В��x$8�
�[s3k�F空�k��֋�4Pu XMn� �B�����ȇ����B��;��$�`�ڂ(�'���G�6�&	X^�<풺R�����[�x�M�sz�1LS�y��x��m��H��������:C�^�Ya��97?������I��p���	��՞�7	u7���t�c��(dĠY �|��K�6���01�X�u�'�~�(l�i`#��\�C��rѸ��D��>-�5[p��VJ�Z|�u�z��O%1M�0�:�ʰ��g�o|��0�lC�8V����d�{50�������boEG����A��?�\���n*M1���I��TE��'��N%?���r�e���ِk]6�Bn�� s@l��+�R��jl�ڦ����IX.���:��T�^N�-9g�n6�E~s_�}
$�h�����b�%�$����vo?_K��^�0�&c�&��qJv��s�;l��p�FT,���h�OIR�Ui^?4���@���X���L���+�X0V���[e�c���Щ|����Ï��u��K�$���b�aw�lw��Y�{��YXW})�M���ٔp��u��KN��� �w���K��$CX�Mϝ7I@�x$I"4�����t������K�V�Fmj�9Z�	�rR>��7 D-���`H$eÍZ�,��]��)�+�t��oZ�l�v�lh?��r�����$��ȷ�qw��<-oRr(x�. ��+W	���ӓ�E��v�1)�v1�>�J��.Ѹ�݆��RO����6�b]AY�,��!ه^�h^�#���Z��>��a�"U!xSo���E���K�ƨR����h��m��nG�ڝ�VB�D�5�����X{��>�X0Ȱ�ّ�5y`	5A�!���y���{ԓP��-1N���BW����c�è�x���߸�B`�6SLs^H.W�`�B��%�K��˹v �6&P3@���16Op*g���v����ke�\�s2�b�A����0z�Z�j���,8�C�I�:=��pk$5�b9�Q���G��W�� ��`��^YJ=^E0���HM�\��S��ZsB؂?�e�Ǚ�c�/x�bTB/8\��8BN�ޟ�~�:Z���63�֥�wLX��_+N����AK(�H�<ņgtعcڡ��l�����*�7J��y�H�Qa����U.;eł2y�����K#��΄�,=���g_�v c�8��M̘�eb-��$D�|���a5�H%�F�)�L�/�W�YC���麍:_N��o͡��HGoV�wT����I��1Ņx�*�kq���J�y�[� ����H�5"(��j\��	~7�#Q���	�{c�]��2o�V1��%)0.�;���]S?�4�uN����:��f�7��L����N*�y���~RH����n��ܑ���Ic��"�6��J�^�{����G3�l@Z0Ě*��}ך�b�{�kJ���jث�v�I |��b���p�l�� Й�y���"��$�(���*R�(�1\��b���v�R�i}`��%iy�U#�ܞ�4�&������9l�Օm�m@��g)ï_��@�i�{/��ч9�~����Y��$�w��_�L��،��B�e�Eb�iֲ�7���jR���R�5{VTXAsع$��ʩ2�=����)���;)�&���ԇ����J<r\a��ȮY������|mhk�'�
�h��{��\�I��/�0C=t��=���2���?��ʠ���R�xIA�����L)\X�?��	�������`�N�W�v.�Qv���a�U�z
P�k�J�4����ر�=���R�D�ӯ�k$8�=d?M�43�sK������C״�ǭ�G`�[T���'(�O>�c�b�go��Ry��r�Hj}�Um�!|��Ґ3La�?h�S��C��s� ��W�4\\q3�
�6i��;c�_�)͗I����P4!�&�P���\]��е���g*H�\7j~&#X�D����F��j��e�A=�+6�{���;�J�JPQ�����iR	�륆�u���1%q�blZj�zG� Buj��E^��.�j��g.����͈/PO,�/?�ӶC�Ȯ�kX-h'}��m�Ǳ��9��4�A��RC�����q�f�G��D�R��6J~2s�+��3)$�$x��o߼����P��\�mTTt�/X@�C�e���ar��}Ê6{��u���Li4�ͩa��%�nbU$'�'S��L3:���_��G���$��.s�V��*�V�S��+� X)�vge���ڎU�����Qov2`?)��:/��)J.�T���Bb�$�e��Z�p洷'�����Lp�'y΍9�j�S���VԈ^���5Q�"-�]���Qkd���;%q?i�'~� �\,Dh����t��LOڳ�N�N�\'�wY�-k��������қS�,o�����"�g7�y����[�v����c�?���ŉR)���i���+����px�����i!_�����x"�vC�iX8���^�SS��ݑ�E�8�bJ����'==����|1?��*�qHS�Ԙ22��ϗ:�U�Rå s�멺h4�Ǐ�_�<��G�Z/ԊF��;U�	\*np��fg����\#��
�I�Ʌ��*/泺����h-C���Ϯ0}�,O6)ܸIF��q�9%>��s�����Wñ���Gщ7��4�!�:��A =�3����Z��25Q,�I6�C����6z��+*�_�s*���\�D���T�A��&�(}h*K��"L���,O��1�� *��v�j"��E]��VF!�7������_)���9[Θ�=R����9?�N��@����BL�������&�R�{���!ǖ�h�9%"�����qC�Y�������=A��R���f�/		I�-䠼i���
f�M�Ք�����s�ɎwEΆ�����#����|c�/����,X��N@1�h��Qp�}V��X��.��3T�#HbW$�;�Ք��AU��*���/�*�V�,M<�^uA3X��̕���H{�@3��v=�:R�����񘎍�g�K�޳�J���\6s΂	.�?P�{���j�����{IȆ�y,�f�8xr��=���a����g����]�~�N���?Lә���A2��kQ����H?Cd�S�F7�K�Ч��U��t���}Ա)\�
w��{1�{�Ͳ��h�;ҙf
�̈́maq?������}�;Z�jq]��L�.��r2Жd����mkՁޡ ������O-x��D�J8�=[���t��>�'��_{� ���x4��K$I���~��sR��G"n�A���:@r_��S��rW�k�=&�F�Ӛ*P
�x��i��� ���2,OGn­m��Up�rw7`8~�6y������l���|*_#b&ֺJψ�.�����	�3��JV��)�Ut��V��F���� ���<�K���F�,�/ށ��~uxH����l,�Lb�8fb�IiJX�A�zӊ]�Uo�YH(��Q.k#�����XtT
���k*g���6�	�����8Q������-�_�t�8�Də��w�T{��V�N��\�ñ۟�6��bW�vf(Ft��S���`l6��	#�m.!R|d��+Ѥ��'��y�]|�ʧ贛A��b]^�/���DU��"������>��}�#�r��ǉ��#�"c齥g�̍z��/���9�~Jfm�M�;Waj��A����mG�S���I-^�D�=�,R����8�'����7H�ۍ�Ё��"p��P���Y��	c�`ӟ�%��0�1`�G��+��2�L�����ȿAj�*B/�����C43�=�y�0��K{[���S3��������-�t�����}�)�P����rx�K��:K�{�%)��i3�F�m|ͣ����u	î��&�5� �uU+��8�V�����/�'��7��6��a
�/x�1f�ǫ�9#��1�����Z�`h��BF!�>���)�T1��`YS?�*�����k�=H����,�/��<S�ȋ�L��k�|RX�l4R�p ��Yk���"�W��!�6�9�{Y+|;H�!4P{����\����>�n*�ø���9�^>��*�56#��fh����k�.`�D,�8�1�s偋��F�,�X2~$V �'�B��>�`�	�FH͎{C�LлǻB�W����C�Y�I@3�Z��6��_�J8��y=�f(�AӺΨ���!����P�C�����E��o��4���'\�y�d�US(X�����������aVڥ��e��a��
��z��iյ��R5��>�J��o�?�< ͎�5W�.�%�U
��\�G�'��\�sճ0[ �h��*�pj��a��u]p�=tj$t�/i�1~���̲�1�������%]�i��z��CV�O�����Yu".�ӿ`O'4��޾��5�"�!
�-��Z��;Y�Q�\aM	0�����V�e���ܨ�XJ2;�V���=�O�y�rN����o0#�~Lq�r<�D���m�L)t� � 3I=��������Z�zu/�o�Ng���K	%�=|z�[(8+� &��6�oy�:�pp{�V`@�h�˶;$E������_�I��?�Fu�H@�,l�A�4�����/Ķ��f��`WV�`�l>8��閉å�(�PM-�1ʈ6ڋ8e;g �����=EfB���v��\���<^��| ��{�Ź+;V���(v�8j���^Id�w��Ue,�%}����;*�͋�lJ�Rx�O�B5b"�'R��SZU\k ҇_w�og�ŭ�LS�ЅJ�w�O/G�˩5m�;�+F̔��;���q�ze_���^ʫ����#I��yqJ6�-��3��{�j�M���� ��0�#p?����eu��s�WB��c�2
�"���ֳs(��p8|��O�f�vʀ�*g��+w��x��*��E��&���#�\
�]�8�����i��/�dD�	!�8���s��2�Y���K��unHO��"�����9��3ֽ+��M4�#i���\�0tԬ�	�\Ԫ�d��ojV�`Cڡ�Ö�{�ᖀ)y�7��g1ݻ)&�c��-�������ʻ��q���I�m
h:�@M�!�֡5R"�GL}�2a�`::�~y���HF���n	���2߱�\Vф�t��^�Aՙ�4.�r����_O���~?ύM��Y�;�m_	�~Pԯ&I�,�"��E2�e�f�dU�{�i�1)bN$:�F7&��t�	ɬ�}��.[�7/Tr.?r���"?�8���z�3�I)n���Q��{-�#�H�E�)w�
bj��ڮ��)Q=S�O�Ȁ#��)��M���d��I�_ (�M?^aGp���;�: /&�(O�A"O�"���B6�iSfs���
�[�m��S.ǹh2"r���П��[
֊x��2��� =���.��,%��1�S�	�7�n�j���{�׀��e�Rq�S�-v��c�'��!��]�0p���Þ�O���N�b�-^��wLo���8��!����;�Z��打����N?�)	��F���z��y���'5X��y�n��/cd�>�WN�Ǥ���F��&��X������]�T�[���F���bRP=�\b@ɺ__k�{�^������,�|�RA�X@�
g�i���wU��q~��nHBnL��UF�^�908x�3�[9�)��V��\F��п��zX�n��[C)nA�*1���2��&�N&�4s�K�L���T��YuC���׀L�[S|��h����)�m����g�� �[iB�0pQn<�K{��.��28���u�"���c�#��*�>#}W<�>]`�A�`�+��I�� �2�8��e�������]
�-k����[b"��%	F�3j��N�k �$G�I����5��g�6���ks��]���s����r�YΤ}�=�hF����|���>w�匋~P�~���p���[���� 7��������"�c���5���K;�� �z@8��1{z�x�7���cq�$/x�B�����\ !ɰ_NE�?Q?Ԛ���·����L�e��#$:{<���
�ݩyV+٦|��x�䊚���b|�&��Q���4�84m �p�8�1���⁡!�L������P���.��7��0�x�.F%�W�8@Ր,8:�O����Ib<��Q�(��r�����w����c�p�d�c�_s��8瓋B�%6�_0K.����U���!n����u�g��;P(`z�V�m�r}��y�Zz�f��#�"�f�*�Ze��E����м�t�e�*���d�-v]�U�h�);Y�@���)�:�ΒJ���y8GEi{�ׇ
��lX�k65��`��T��K��>ƴ�J�s_n^:�qy�	_,� ��5���o�3^,oB��bTKBD4$�9�>{󋥸�����r�)������2D��c䘞f�V����O	�ݴƠE
����P�����KQ���_y�,t�����J�����i)-e�E��4w}3Y�BZ��#���д�|�HT��Q���0���!�-e��\��;@�s�$Q��	���7/��23�}��<�!K��7�~CjuI"���h���5!���-B
U��+gPw*�i��z 4�ew�;��VV� ����'gUuZ���4�n���䘓p��DXמٗF��<vF��Mغ��qי��j8���6�f3u�7�'��(����.dܨ��4��d��}�����Aې�O|\�2�L�pe�Va�X� !��#ݛ�M�1�j�=�o��C�/� ;a8T˨��Tr���H�J�:��e[��"��]�ZJM��~g��z6iO������
������������������IŔk͈>��;@z4 �%���>�1���j�x�w҅���{X���v�|��%\�/9
H[��JCif׬!��.���Ҽ����;���O�˫��,�i��*��-+���ԩ͎HP܊���!��6����9��b]=�`�=�͵
�&��N��u+=�3k�WV�1T):�=��N��8Q��:�
?���sbg���F�d��8(:�)����b�s�C83�9Ӫ��yO�����?9v�6�&�נt_Y�ɇv�Q���imc\@1#�A_K~?VLt_�i˕�b�h��Zgh�����2���W�2-[��hbR��O��w[�q7�.���90���^��"�N�����:g���'�d؉�Z���'�Ǵ�^��u�'�g*�3w{z-��yu9�lq��i�E�cޮ:���hf]���!u�8O�zwv�^Pyed� ��XE_1�N��-�Mjh^]��"T��A�5�:�<�����∥� �P�Xw� =dm���Y����p�F+q8�L
a�o�C>�N�XB< �c��j���H$i�i��A�1�(Y��*��nU��J楘���7�a"y����j�_=ҹ����)���˼n@�3S�l�����^+�co��K�_Q���x~.�!��{�K~י1m����^ed�q��E�L�w�"�]�.u�����e�ٶ�N"�=�<�5+���7��{Yt*	�_+�S�j�x�����G��n�%���tDˏ��ŉ����|k=N�^��<�laR��^�o�h�7�z�O����9?«A�;��-Zlk�u�l5���r�]�|H|+5?C�������Uۈ�ca�� ;��+��W���&\]B�LC�H�9F���r����֧1	��4�Q�Py_E&���5J葁��Lb��|f4ٮ��8�G�K8"n����_O�:�}l��ߺ_;���>G��NP&H��g'����ҋ�.�K��j�4�S��;��8���t�����nY;f�욣'���q����6� ���f�_����>ι�GG���	3���«��1K��p>�(b�Ď�����������lIC��v@%���
5C�L8�q�����n'6��Vv��k�������P����6�ؖt��J�#u�R�m�����X3����-��5��1n6F�1��렼S�R ��P���B�p�b`��/�wl��F��쓟q��E��V.x}_b]�@]mhBR�̒��)�UK�nځ�������F��x�B0�`, j�*o���r\_h�usI�3����]ո�����}�;�ֵ���y*�33Z�ơ�(#�ɑ�c��
#n��5��E�r������3�
vJ��6�>Ê09��74�Ft7]�C�������v8om�'/���R���1�}��Wu?����y������[!��u�+x�B�x3V
+Ɍ!҄Q%���Pg�>�0���+�gƕFV����8�fr�4Xf��]R�\[��t��k�<(I��8��������Z8��G�џ�&q!}\�[�#��@�fC�u.�(�U�)�	y��!"�*��>��Y���z,`@ʩˑ���$M}��E���)s#o/ ˏ�s�KS,Z#F�%�p�+�i���֛���36l�U�RS͟��U���G�?�`j���0\^c���2{�@\)4婓A�S40��_GqO��%>v<G�:�O���5^Df9&)��
p���oJ�����`$���U�9|�Ś8���%�ە����7���9!�+E��3>
-���0ȝeB�ny�m'��UaOɆ������> m{i�o��;����Kb�c�f��x5�`%�GŇu����8Z��J~��s���↎La���&���0�%|aqnWǄ�K�q�,�Z�G�x�SkzE�	�΄��~�q�5��I����=�TqL\��!�Gs����nϲ�(�C�ܶ��
xw�x�bW�=���p���9f�x���#��^ٖނ9{{��f^�4��B(}��n�s1_�r��F���J垲w�=u���=�E� �����M9�2����x�7?��9���+cP]0E��|"���ɮ��\�����`?�>`���A1�%]-�@>�K�BZ:[�6n�9O��M�V�n�%P&8f�J�?�*{�Kw[���u�à�z};�\�`k�*s�P���jO������f7�	��	�������U,6�o���']R�3��s��}@�,�ޘ-ٖ�E�|�ǠYӦY.��[6��<&��I�w�W�omsX�����+9�A&�$�YE�J�-ѩH"*3��c�	و���=Ϧ�����6�vL�=郺�R���/_�;o�ͰΔ��n�Haa��h�.@c�rY���
��&�8z����JVD�D}�~� ��`=���7��D���1���T+�;��=y���@i[��? �t�|�c��}$�8��A�ĝ@
�E2^�,���sX[Z�J�<�B�6���h��;[����g�g�-XS*�$��8'tQ-::�xSɃ��&-�T�ݱM����̺�I�/I��n�͎��0ד�u�:���<�[��Z�&�#�;և��M-�1�
���	������U�|攠��``�x�V-@s�h��&.t}O1>w}�_���he7W/=�d�*�N�2AH6�5O��ΊK� Y�󆫖W��<C9V+�0�N%7�"�<���6ea��V;3�ٿVJ<�:��,6@�u�K���#��������;!>��5��-`F���jDS'�J��v�T>3{L����L���<�l�oh�K��un	��X��$,J 8k�U�:����nT���x�L��孽�r=f)E�G�A��i&��GH���~IWU�7b�@�z*��\��z��c`6�
O�rD���/�/[P������qN��q#ԉ^^!_�8}K����_umI�֫>S��.�w�ɅU�����+��3r�[�;,���E��R�}��M�>����{�$���h]w�{]��:O����=�T푄ɚ.τ���7�2��o���7�a=k�1i�ß���p�>�];4|"h&��vy1ˡ���M�Uє?G��{ZW7$���s��-�D:=�wp�zIF]�<�9�F'��-����))#����wDt�~վ���֯j* nh���ׇ��5���yʲ�2Z+'^��4��E�LLL��E�"d��B->�"�≯Y�i%$�V4�ļ4��LJm��=D���;x�?��� �,$��W.o�Ւ� �'�x_��(=6�Go��y�ð���#�t{S�`Ѝ8��� ��lb���Ţ�d�m�~B,�EY�H��Sũ+���9������:�5_���j�g�d㘺A({K'���T��6�i8���>�,��wϏ!#�%��֦�ɫG���+�+��C�H�	���s��7\���^�L�%M}�ݕ�.D�@6������=/U��'P��Eڂ(�����]����"U�mc�"��܂�oB�!�$�+�M�'/O�m�ت��80��qYT~�;������}ޗ1�A(wI['47��!�H%�[|��o�~�3�7��xiY=�v��t�n��;Xt��уJ��SRJ-=��x���k�W�:56�L㧮V�h,W�iƁo\�T�|S*��~~A���Fo�7R����Ñ ���nQ9H5����cR'���p�x�]N����]v�������>������q��s�_�	���h�72q��O�%�.As�7��U���$�~��4�j�Fpw��1�@�^��Y�}G�ql_����|���8w��ӣ�(z��T��.]���̎�g��s��fQ{�����D~Y@��;�j� ����U0P_�HR�x)��A����&)�qMY���wM�G��K��A���l�<"�7P�EI� ��R�'���������#���S6Y��<�\���th�e�L1���;�k$��^�!3.�6�*�$���0M"݉J��,����0Y��l�T�tXZ�c(05(N��rJ%�v�����[@�irK�����X0�E[E�(l]���̫O���va+�s��aCs���?}j�ڀ5��<XR��U�3E�@�
����Y�`��o�$~��O�;�Qq�)�rKљ)K���7�C����,����f�u�>���[�&��,S����l	Yp�M3x��j����8�5��'E�I��Jv@н�B'�+��,�O*���"=��t�0hC�v�ؔ�=:�l�1�� �0Ƒ��
�o�V[5.0�׼�P�>+��߻O�m~�j����V�������N�*ރ�$fGo�j+��N 
��K5���c��M�Y���Q
��m��3f���"�.�.w�ʤfvH~g���@����Y�r�;�W�nc�\��d�Ňզ)٫pBs֭�U��bd�o�Zv������/l��Q�fS5�?��Z���j����UV�{g��z�mOĽ�@�Md-)@��Y�w����jT逥ʱ��w�"A-��&�J�Yg�Tv��
���N�
j���X�N�ؙ��7~h;��E]H�X����KМ.'T\��s���Z�'^˱�%*j�}>�SY۾���w�Ja���MDt�����F��D���Uv��o���k {���1L�;������r���� 6KV/j�����TI�e��]��E}랫�X)1�̰�M�dYH~B�K��{<f)~DK����h�Uk��&{��_^�8M�|5u#ib�v��Ƌ��_R�zIѫ\��;����(��+�_#�+��6e�'.x�O(��V$���ڭ#�۝�8fa��qH�����&�dXR^��F7e,(x	�d�����1a^��}]�1�d)��Sz�u���~�c=��?�x��᷽��e�"��t^�����/�ʨ���BH��0�EhiU�7_3O918��1��l��/,R�;S�	�H��HcAP�0_$�BKwx���	�UKȤ}b���Xr����Q�j�Sh�h!�V]�w��o�W�x�{������#5_ͼ���3(���8I�k�'�~(L԰�2�_�sX�	��?axT�$��6��x�6=�鿠A*t���V���Ҙ}eYBV��Q��y���{ZSZ���_H��p����`�+���J>�+�X��qˀ?�� {)��ثU_e�N�S�.��2AKo+�C� o�[�u,��;1'Ŀ����EL�M���xGٝ���vC�m��o�X��P�s�c�t�򔵉Jm	����(jI�����su��٘��ǽt;j�&���/{
Q��w���g���*#Wͳ��[�)~7��-2w(��oJg^C�D��P�%��Q�Vk���c:D_:K8��#��!�t�Q���e�όR�~k�ǽ�.~޲��� �PYx#����7v�P;���ڑ�ȥf����!�襹�Z+�
���"f�#o�X���U���s�&o���/�vPt杆re�p���Lu��Ph�@�č ����U�G�g���*����`6x�9�R�O�ǃ,*��\7
�:�d�0�$4W&��6�UZ�M�c����u��O��'���6g�����m	V
^#VJ�
�h��$���<|���5���|v��;�^,#�wݤ��~���O?��|��q�M>4?,��5�0�.[6����,}��#	Y��Q1�9��27���-��HZi�D�h�ԯ����������3g�����I�#My���������X�w`�>��9i�c=`&犧��o=�}H:��jH:��(D��p�Li"^���]-�+(���M �b�[TJ���h�1��������a��j�аR&��)l��~���nM����Γ%����8I�HI�#�d��^V�7{I��B�����OB�^��GӇ&�/񉶫N�_�i�?�Ы@٘������v�`~;����1�R��|��4�����}0�Ң��y�A"/.�)��q�.���֡���~�	��b0v�8}��C^t���\���('TA;�Rj�M��\�I�V��= J�(E�:~	�R���鈙v2iW�z\�Vھ�-,�4��D�eО�/���7�VY��6δQQ��ol��#���1M����C�>���9\�<b�b�(�D����0!�m���L-v�x���cjs 58���wLs�z�n!7"�D��L��i���T�ǋ'�dGT�@� t�!���-�Vo=9T�(J�J\��[�#,`���9<n��4�����R&Hw�B,1�f���0=Wv�{&�Ɍx#���<���]���)�&�B�@ �B��%��}sw� ��G<����k��h�Q�ֽ�[�k��d�;����W�x�c��98a�V�-L?�m�J�����v�x����v���͈/��ǭ�6�{'��m�|w����cC�d�ĉ��?�>����c��3��f/�?l�0�aI�Mghy�R�ZTN!���ߋ�]�*S����l�{SCc��M��ljnl3��R��K��.�p�����(�?��:@F�> ���˟g��>Vv-�.��ǖ�����?<%�'�P���H��6�x�	� P�#�.[������dm��6����-e8sT�,��R�V)��|p�t���)�/O�c
��y<��S�hy���ch��sװ��҅L��ԯc�� H>y,&^z�E#�vqI���S�+�Z��)g��h�b��ں�Z+�[a��TLNZ�f>��e"LI�[�^���޹���靄��q���
N�J�t��Θ0�A��Uu 8\!���wx[L����ew��i�X��u�%Prթ����Z.�TZ��?�����fc���NRX�s!(�5*����͛�¡�C�#k�8[f��S�����7j�t���� �}�
b`�@�ea���Ec��Q�U�z-*c�VRm7ۓ$k�d��������=������/"(��W���K?s+W~GZk&��+���.�HTƎD�K�J}L��zC]-_��e�
w���jK\J�)���s�����aUjT�nq�0��#)۳l�Y�kt~��0�m����}�l�oc/ͫ�0�2�(UR��������ٸ�_��p���	�f�|դ��.?��Q�O�#C�H]�3
����S̤T��)�x<�oȅ�@����L�d����ǐ2��;H�=r��@r�[xW�5�wm��[��t� �V��<�ϓ���oٱ#��y@�Y��#<�xPI�g�2���\��"�2�o�\�n�܄�<��`�	��8M
��<���FI�f�N����&"�`�O!L�⪇l����LV��1�-����p��?=٨���+FW4�X#J�:�k��Y~Y�x&��wK'�#/x�M���P�[�3�ǜ�hx_t[��(�ݪ��ִ	�4�ҼN39=�=t�x2�����h��7a�W�C�\ޠ��k��*!"����+���6���!"��Z-��e� �=�'�E(����#���)��Rs��_��gM=�@`�ii{����fp��b3 1��s�k��@��
ib`��Ȑ�"��bL5��8%lr����3l>g'Uj�#R���1��˖�x�����B8��΁��Pz!�j�j�B�{⩳iF/-�6u���Ux�1�xC<ʵEIc �8�4Qh��rٖ��xO4�@E�^E�r�-�L��zX��OC�����
Lʤ1��2.�Q��2��,���=%�S�kᤋHq��.��`kt>�s�?C��xZ^���{�W�Z�Mq����q�ԢǑ�'�^>}O���C��s���^[H����>:�k}� a%�^�.�cO� ��w�'�<�~����1	潰�=*�?�׭�J79��?(���@��%��w�Ԯ��9����S��ӧZD�a����!�o[R�4pq*��5&Fu3�d���^*Ɛ|-����x뵩�:5}���ѻ���'-(��ƒ���%�s�p�4�5�X hJcq�\�>��y.C*�����&��D��զ��W��B�
}o�mQ�"�����!k��H8�NyY-te���0x$���T�cs�3���� �ب~_31���y
ߟHi�y�|Jb��_
�x�����[��e+� �٬k�4�idY�������җ�5UhJ �� ��$��Uf8��b���u�2��%jiGV��\c�멝��[P�R,�μ���6����Oߠ
�
���� gv�v��Lp�L&��J�f��!t>�.I������H�%��)�l+|�M�y����(�Z	�z!/.��p���mr�t�ݬ���46�?x_�k3��4�߾��w��ϭ��r�k�a��fK���/��!8��zs'H��٩x���������?g<=XB��B�1&��+�6+������sG0��Z���GU���Ɉ$D��,�J�#m�T���7!���1mR���:�Nc�<�O�2����	h>Gn5�V��g��Rsɶ/}����j���D�+���t��w� �/;K�9w�u������6b��kN��$��;_s�lka�O�n��4J��o�PA*�����R����TplW�5WExY�E���Yk��8Z��0��ע˴S��Ҳ6���*��¤���4�*�{��$�܋_���L!���� �)G�%Wj�`�&�T {h#�˒��巏8�{?���B��G����m@�\[K	ӟJ��_�kꎾ���C��xiϻ��ȩ-5U�N|�R��vr�c4وK�U���F]�4�����.K޹yX}	��յ�w��(���i޼ܢ�N�m֬��w�#�ܪ��;�2E8IT
	�Y�Fd{ff�z��%��̞��Q�ЕXUoX-scn�׎���*3���<�1��*E�Uum�'o�.v˚�:vZdo\�n�I�n���H������|;�1�.H~�j��t�����bf��a���Bj���ۈ�#��b���B�3<R�a�����O��靗�3�_���]=�x�3=+�g0]���=_>�}���Lb9�]üH��Y�f���c���U��0v�.(���ˤ�l�/Y�?�c��WJ���`q���:e�߳���������C��V�E<ܵ�Z,f�f��t�/�:410!A�28B �BKgؼ��:������_���T�|<�C�^GJ����ĝ_�݆UJs�!s�K�R�<����]��j	e�Y��,�0�Y�& �[��rv7�=eQ�j�Fb~���ҩק��5�3r}ho5�/��";ڬf-��-Q��+���AM�����%�������N/-ۘ$�@�l5ʁy�VTIQ���Zz�̌�ۋ�����j�9?�ȝ����&��֥/�S�ND7��
/U%8�`�;������w�8�t��t��7����(������q��-�˗V�CY�e3���EwB��v�j�J�#�"M�J�9h��L��i��U�5��e��
�í}C��#Z�!8��5��
#(['r`�	e�5i�2�����I��5��&Vp=�ÜO>xVʴ� S�@����ӘE+��reF�F�ʣ`�A��B�����"����k����k�I�/���
�]���sh���b~(��d[i�	I�_�#{���q���?����ᆛx�
Np��)I1���z�oW�H͇3,uC��舱�γlCU���,�Σ<�3��1H��`��,��s4�r�wu}̰�1:���<R�o��M�F.s뜥��	����|���ئ�j��`d���0\�j�/+Q�tyH����5��A:	���)\�i҂v�D &h�D����q�/��b�J���pU����8@��3�5�[��%tJQHl��g���g��7t��Q����L�b�&e?D ;1Բ����7�0��J�dt1��P'�����y8t�����p�^�Q\��}/���C��8����l��?9�8L��=�)9�2�.}�M��Gۙ�ŋ�ɉ`C4�V+3&e@]@�#+H���D� ?��ɢ�g~�����ĩ���͇���u�����E�K�i��[^�u�5������@��*͸���"/��|����	��[fD�a_FZ%_q����}4�4���/�bfAi
1J� ���u��P[���4��d�C�@��=â&ۗ���1F ����A�j������ނe��D�l\}l���H2��_a�,	5}���u��!'04(����ߎ=�S����3��Tv#���"��nU$ˢrW� "�m�Ucg��Ȁ���f#|� oV��n&�P�9�V��W��EkH*޻ޚB�}�%���Qk�
���������;u{"��܈���l\[��m���[,�����z�l�@�8�t'�� ��_�|���}S�O��鶦z-�s:ԣ�w� ��%."i(��Ͱv�]���y����]r_�c3�K���}��(��E��ǜ�s4��O�s^Q��4�/�A�*I~�W<[Û .�fׂ�l�*(�s�I���fL�x{��s���12��K�r& �,/�[y�;����u<4A��i� �H�AE�T�?j�Ѳ"�أ���#���ᕪ����E�*C�����~�Z�ȏ�p\iSe���1˹�P�u��Cz�0��q�P+@T�(c��q@�"��>�&��'�Z+Ȕ�uVL�d���g��s�#�6Uʛ:�l��!+�w3�>���� �&�G^�$�tJ�cՃA���D��j��	��i�$.�:���ڷ�y� ���Z��c�P���g�æ�_��&�/�>[���������`G��1�ёP��_F?m���f|D���my=8c?�����.0��J��d�Z�.&��bY�,��XY����Y+�	�h���>"]�g�-y�6[D~�8��aU<\}t?�&z�&ע��Y+��~b��/�Tz�

(��j!�xB���ŋ>�F�؆7+;x���� dd��tP�-W�E��,ݩ
��Fr��Y�Wn��蘗�,b���3�
	%
#�����j��k���W�V�d|?A�a��Q�B2�3�I�S���%�F�)���:;Ka̯��i�&��A�7�4�P��"����ɉ�f����K��A�9���������n�#���D�=Yr�&���s�+�p����S�� �R��-�b�a�A['�7�Ap�n־S�{V\��b�_�I'g�qS�Ե�����v���tS��{���h��5Ȕ�tًa轅��N�	��z�c����F5��!*i^L�@����h7�Z�&�9<�G^�"SM�Y�^F��\�%A�9^�ר�0%!i�;f��k.3ګ��t���r-�_�n�җ�%�Ed�lu�R�����e��/�J��L�V�A1�)����q���$lWv��C�%�)H���m��,6d���:QD�����(���dGeB��4�Č�{$�v��-�� ��"��?���rOR����<�%}�����Ґ\T�YdF�ȶL�_@>�;�J��|�Yb��uNㆈ��za V5K��\ڡ��ؑ�����K=��(7�(�h�g�o��7�����َ1r`��m���XL<�(��Z�VT�͑�*H��)\v����~P���N�1<�Ń��������':�g�ڃ�$5^�mSe�K���5�BW[�M@�~��O+o��5� ��|��4�� �A�mr����0}����%�Ū��GI������S጖K�D�9y����ybB<7�[�'�y�;��mJP�S�35��_�'��,i�j��rf�d�R��Υ�/���	lh4`� S3�a�]�eh;.,(^�<�� Ǥ'e��pgߨP*�����(����D�i�j�A�s�k�S�mp;$�W7>�����cS�h������ڟ�i�}� V������z�V��I�xf�z���Y�xp�NQ�p��Lr�H�����&<�ft!.;����Ԏ��-_��]3�D������B�� e�#T��N##!Pص]UkcWgA�|��Nͨ�|�U��ѫى�r��b�����p��S�"|� �2��"|��M��Q������蠐D��aM���#�g"ɼ�W�>.A�5�kw%��/������.�g,6n#F��0���]��h&lN�6��n��M+$�9N@����` 	��`P�T�n~	΄�����X��d9����Va����mJ�g����%׷a��
_@ �����.��=�Q��$}���˲�U�sm�[�(]UCBl	�Gz}��E���D䮶�w��q�i�"b����k�d�YY����}�pC���ȷ;����"��f�u��aK�Ќ$l̒���s}gM �4eK>a�M~�)-t��B����¯9�L��,�f��֡�n�<Q��A�^�V�P�KWF2(�*�,��q���O�y����Z��p��#ۨ����7>O�Q�;6�>,�wg��ꥮY�6�b7��]x5�+>���T�:�kD�M��2���o����\ޖ�E�����q@���oIqB>j־�F節�I���2�9+�u܄�TŹ���>-2��/.Qq�?
۾<����qTV����!�"���.�)��A"XUs�IP�a��XD}�ܶ�aǌ)ٺ�Nv���%�v�$��	&���RAl��<�2]㖞��VQ��]wp�+8}����xD�(XR�x�lJl�:+A}&G�����Qn��֬��<!�m�~P-���z>�;CD���P5����W\Y�O��p!�?�s�X���(�@���dR��f}�x�|�.fxM"ӉC+7�A,
� �8�,sV��}�(G�>
 ,�����;�f�1hag�`9�Q]��|�z!��!��'�'�JX��16�j��I�y�����"Х���S����di�w�2:��CH��>���,�����)e��Қ˧�0ײAJ�V 3��$L��8�^{�����Ủ乲R��Q�,V���*�J���X�:�������[��L�N�˕L�)?|-������$p���.�؏�!U������W���K=�s`:���~ݟ�����>���S���N=?�Z6������&W�y�E7)a0&t'��-`�'1hS�A3����"�&3ߡj� b{��#Qp��<,�-�G��+w[�>�~g��N�)�c���fZ߻���MZ��c8�j��������5j�:��묛!y�
7<T�!.�,��T~�&C�Ma;?<�	���4M<���:�q[���cvu����:��V@@�t%ˆ��bt�J�r�?��F�)��]�^̃�+���|$).ɹ+lOb�l��������`�qi��%5��ҝ�1IS��u��'��H�=������/�����V/g�w�aD[܊���e �nŦ��*�x�j\����?���=V8�c��l"���5X|7�GY��>�<��?,�h�|w�T'��2g���$�;�if���5]t�<+~�m�X�kp��Qt5R(�Ǽ�\*)B�.���.�A�Z}+�u5/  c=��ŁӪ�D�.@s'\����qê��%,���7i�%��ߖ����59�����:��SY�*;�^����y���ۉg�}�����
��������Ӟv<� ��5P,d)�9$��l�MH8���r�5�5U�]�f����(�/�X_H��b=x�^�v�ؚ10_�5��<h�qG�'Cn��> �;�w�C7�\���dMhJG�x��\��{z4&qF�jl4�� ��J
��|��h�����& |�3�W��G(���l�01:R�u����X`PP�o���0W�j����'UA?4D8�XG��b���P��v�g)�\�Z[lq>M��Fz�k���Ӧ:v(��W����^�X/ɖ�)�n2�H�l|])��1"���]�%�H�޶� a<�jVI����U���j��t�_�r�4N[�4��M��͛[���ѓ�8��P&�w=���s��
,�w�͝�<��Z{�IYԀh��9w��S�o�AJ!r�J��V���{�QQ��ӿ$\����`�8��!.
)G&�Z�����?�-�?4����4
���VS%���7����5��(:,�S(`6Z!�L���BPZ��ޝ��?��=<�������I�͊���;��s�����^Λ4�����0�0R3vX���l�4�ΕJ���P��E��^�I'�󅢘��`������%�_pK7�(=L�/:�p��2�4� }AP�t�uG��X
��ɊX���>�Y�~v��6lڹ�"�Z��;��+��LqڔvAy���$G�>��N~�^�O�Ov+V<c�Ӭeф�������ī���{+Q�9���؊!�a�5`4~�M���������X�u"ʫ��H�)kj��Xk��j~�q
��r^L�?�j�u�q6:���_>����/�o$ U|����~2����OQ�q��줘��`�N^�������m���&GӋ����2Mkܲ''��fi��q�$9���$黗�.�fQ��:�9��6�sP�U����:ޱ������`=u��h��`���Z����ڑ6n$�'N�}��P�E��]t7��c�=��:�}xiЧ�RM����+��.^L������ܚ��ՃCL�3Ƥ�k�b�z��D-M'Ɵ������n�������Xȋ��j8�>Q�)�A<2*���~�T[�BgO�FXa[+��2K������w�@J���?E@��ay���+���&��?���9�\n`�v��B{��̇:�A�C;��hO���YյD�p��{� ��Y�sx>���%�a�e�u�E{��	����y� 㳢d��R�S?��d�2���3��ß8�1�9J������J����>��7\?U�D5�S�7�7o�|S<��j��/�5�[�������B}q5���a˜��/��HLv4��蹰m#~ĝoA�q7fI���H���ۖ��]���S����<h�s�W���**?f]I)}� �o�CՋ3\T���++�CL@�6�kh��5�'J�n�nas�4�������g��ߊ��@ߛ|Z��|�ň�'���%���gՀ\��6!�r`��aiB쾁 �{1sa+Y�A ����kWf?3 3�zNMz_������N$qY�~A�)i��z�-I�/�;N2���J���Q��3><�ß��M\7*q�v� �j�{�ӽג~2N�x��]�Y�<�t�B>�$���Z.7f1�y}8ڃ��J���J}]�"���W�o�*6l
�˜~����M���K*߿ݯ.���F�N�L9�={W���arג�e�;����g���d������i�}�(k��#����d\N��O�+o2��@+'@���x>d���yn'?[9#�U�,��/��l�f��ȵ7���< ~�����\*���$gg��;g{$�T
�l�F,U��m�J�9#�O��*]� ������h�U����C��{6��{Q�Q�v�s���YkkW���6�@�ᕥ]Q�
&�T����W~z )�IZ��ha������ۛ��J0b�?g��ȏَ]]�6�>k�=�-Xz�8��(wY�;���3�A|��RC�fG�rz4]yv(�%�������"���_��	N�~��I3\��?�l�[��6M���R�5Ş=�-�BGx��._�;&���t[��C��F�	d�y�%q:y�{�KKO��׸�_��QKoh+�����b��!3�������BϞU
��|앢�Q����D��A����h��v�U�ێ'*������܏I�F��4SF������R�
��oQ�{E�$�h�k)�ٳf�k-�.����gۅ�S#�'���z��-�h�/�{��܂>ʎ����S�XVH�������{ӗu����-�&_ѓU����qp�mCRy'��S�'Q)fNrf������D�Y�W����~0�QK���G���Dd�I<���ۭY�t�� DJ�ƞn'���N?'�<Xl.�N���I��*00Q's]�bæ�7l�])-�!o���
H�
�{&S%l}D��t��p�:��I��;�[�^N.^@�=�<Ϡ!�Y��3��g�֏{�H�`ab��g�;b$�*v[�UqC��)���_���#
��\8%��a��ýu<�	_�.ƵF14�ץ���|�(ӊ�D�'��j��n����]��Z_]oNd�'�5�e�6���^< E��j��ǥL�w� �Y��+�;���P�u�*��zIs��IT���}ap���%ؤ�*����q{W��e/�î��\��d*��lo�@�M�e�����%R�5Y@�U�B;�D�c�MvN���IʫW;+�MyZ���g��>���+��O������-<�N���#c��f�`ol����D��&��L����#��7/v�����&�+�j������� 3��v)j<�)D�>UU���Nc�e�ֈ�QRx��D˺[A�1ΉO���=� @A ���ײk�� �?I	耤Ja�#1BC�S	�p��������V�g��"`|�碉���'����I6D��/��ޒ�<�G���
��r���'h�d�_�V�r�u�v=�K�YTӟ�?i���w(�1����=�r��xV�h�S5g���Ht��.�4!|O�.��A�����)t+�<pz�Qh�D����a��O��:"fך�Y�zE�B�ݜ�^@G�?��P+���C���w(�<,>�7���+[���^�Ԋ������A��9��8�a��9��H���^��gC�O�+^���;�N����cT����تa|��u+��Ψw��fK�:JBYמ_��74@��c����U��!��;kHL�Q���bw� �'
g�E��D��E��������`���#w�/�=w�!�w`��������
b��b�>�D�J�g�zJ�4�z+���8t��	�����GƂ��)D��i�ٞ>~ޓ��'*���r�4NJ �HU�6����NKi��"c�Ü,D�*'��8��x���^�W��T%��H�͛�Q��d���� O�#���0���I�C8"	��>�+G�����)�v{FK�/R�������K212�<��?���PWq�Б�Նo=R�U��F:"j�R@��9z)]�B�����t�j�5v�
_�D����^%�݌�M��wl��G4��~k��w��,w�}�9��Ҝ�[l�g�\�A#�\`�U�*"��/�,�4b��h@75[8�Q�H�j��p,��~�f�vx���VN}M�\Õ�1%��ZkH���1Y� .�>M���>�{w�F��Ӽܢ��G��n5�U���Lt������bgַ��.�m�^�ϡ�MaB�$�G���6C��U����nbH��=�CD��惤���{��T�kd�8Q>s�^��� 0��Vf���dgqn�xtA��V�����ס��Ǳgkм��[�ki��$�+��Ͽ)N���A[�ڤ���_{��U��ĵZ1O�x8%���+�9c~�VC�ҿ᪕� I���I��/Hf�o�p��E͆9���B��B������L��3ZK1o�?�0eSt=1�$���>�8��{e\a&m��qj�zV�Ɲ�*8є��˅2X%�x�Ht�U%�O�̵��n�Z�ft��/�X�����tnH1j��4���XN۫%��Ǧ(|e�~�|Q���]ô���Y�fy�����f.{��a�:s8)Yw��^�+��D&n�?�q�t����Tv�f�}U0�����S��mKy�s�
�N��CZ��T��W��^B GS�	PMeF3�ݽ <ރ~m�mr0�������u�.)$�k��­��?ad5�{/��K��W
Ո�}6��|��{��筳���j7b��	�|��ķ,PP\�:�et�ˈ4j,�,O�4m" ����7����V���nV�͈��+R
���?<	�.������J�YM	�_� 35.�9gc�9+�����>f8�L���0���F�i~_��x��8�l�݌�"�-�@8�ф�7��4}��&Zf��� �e�_�l���	@p
9�j
�[Qo�b K�t^x���E !2J9�w�i��(�$yZk>��B��&�W��D��	�����r��7R@� ?�]P��u��tVz�=��5��\��A���/�z�����]�����}�,�;���jh��C�O�Ka�����`��gTD����-nw��C�s����TĞ�)�0��<��^��=�P-�帑y����ƫ{���-�y2�*�|��5?]�����z��|�Eۍ����{Z��_��e��:�{o|���|}$�Z>��F�5�(S�;޲ �����1/'6:v�C�#j�$�~N�X[�6�E�ZɀG�V�{Li`����@;~cZd��Ȉ��[��G�.�@&{F��k�����s��9Q��ܨ�O��V"�ߴ��`���:(��{
1R	|���L����5�h���u&1�a
#2�Mk�K�ОOs:�.
�T��؃^-:f��(,K���5�X{��舣�36\Ύ9!��^��8��&�q{u�]�$0�err�
���٥�
i������tn��-k�3-J��ۯחݫc W-4I�wt���� �z*�qs,�pb��c����e7�7�CD{�|q�z�gЉ��s��9:������m/i���$V_򘪭�H"!�@u���������Ķ������_D �q~߽���c?�M��jQӞ۔Hz��<z�N�Vm6p��2Ha�A2��iʱ�8�k��X�{1�T�BV�� ����σ��S	#�c���.sʋ2�g�ϸ<�u��p��q_��Ԇ���pU�mh��XR�H��܄�2���q�Hǣ^t��*��sH�L�q|.'M�ɩ�C	*�rK�v%F�g�ԭd4�u�<�E�)QK���
�0�R��s�o�	����lg��(/
b���t[���;�Qj�w=>��y�3��k���俞��Ɂ�H�|�Ӓ?�SxY�Nd (��s�BT���R}�v���"��Ⴜw�F��c+����^++��C�΅�C �������Hww���/�5�e��ٹ����b?@�C��E*��jL?�w�n;�o@ruf�k��:P���L751�J��ׯz��r�P�T�Y�W(�[L��-��� ̻HУ�,���u��q��'�W�v��L�qρD�(���n��$SB�k�����7��5�}#Q�-�p׃�������p�Ǐa��S���i��^�Gik��ɮ�d߄wd:��������
c��>(�*
����8��zɐ!u�2vF��d!F�."*��qk�`.��"՜��DrZ���RӘFͳx>��x�����S��3wӣwy6�/�Lh�Acf?�=�s������i#
T从�񟈀\T�vu3��Yu��
�Z�?�����@���_�)mm�e�+��Lck�(�]Lc����U��_�K<��Rf���d���&ݭ����2C�*�G^�U!G���y��I�F�6n<-��ʃ�ރw�6#*�*iG�B�쑰��~�n/������Ɗ��81�М�n��q_�oq��oO:z[���P���B��dt�'ڟ��崴oT������\ �_�S+�t��sCC�'>�J`;U�`b��(0'>z��⁘|��F�!�)���Qg���r%�?K��.��?��
��r�2�q�"`D��V׌�Qu`	Y894A���F���\���t@Z�~��$ҷ�:�C�Aa\��[ҴS� c�^�l(�ɫ��є�q�k��N�GڥG;��!�/�2~Mjʖ�#��f�Q����A\����|�*H�Aއv�$�Ggz��s�;;RA�1�ckk�#� :� �A�[nΆU�굷� 9��b��D�t5�I�U�JIyp&?��1*o��b  �z�D��)G�*��
��U0tI#��;�ڟZ�|�z�U[.@�SV׀J7���k��x���u�MP�d����n���o#괪�n���~O���F{���%�^~�Dd�������pq�h�9*F	���V?�1�q�����x�bht�f��"�y`�a-/yg��`���B8I�+�8��S`.E�\��1	?#��r�1@˕y~h���t�ˇ�V�xX�Ӏ��d��X7�PN�l᙭6��w?�r�X@�)��+k!���u��S�ץ!���)������1��iO%�A�0���ԭ�c»m4K��K�a:ÝD�Y^�Z�l�?f\��@Dϕ��Ɠp�TW]teq-œs�͂T�N�����a�����v8�$��V�$tË��+�u�ƽ/1�)
�K��YOl>�	\�q�������3�c�#�����oyvJ�څE�r�M�&1�ڨ�e�oB5P�l���!������Y,Mb� �����w�`��S�����c��(ޡ\�^�)5u@�)�{ȣV���i_><!X_��f�y�m�>���/2�����"AB�҂ĽlJ"G�3�ɴ�h�Ϭ��O��A d?C��D!T};�(	�ގt�ހ�Gx�(3��qG���4 x�Uh� �JCދڳ��XJ�3^��Σ�0n��|��u�����t�)v��g�'i���K- c+�^�JcI7�0JW�t�����&�_�a�F��DS���`GDC��NVc��C���9�y�"oQ�.��\f�B>YP�&�/77�r��?��~����w��q�,���;�!����\��E)��9���x:{�P�p�S0&�*�P����i�kNh���E���)���:�V�S%�9QN���o PwO��*��L$��L�.F���x�0+Y�ض*�~Z����$��LK���z.O�'�sJ�ɺw�u�7��? �T=��9��-}��>m��6���^c���L4��6�ۦ�+%භ�"�wU��|1S:(#s��ko��j �P�>��E,@���kFCv�W�T�<<\h�̜ջl�T� ��r�P��(�]�5@4�SYX(�s�( ��4�w�Lި���*.�n���^-t6�ߧ=fz��k�DF��}���4<C�y1wxf�;�_���k�.�>F�,���48D$�����2��Ep��n�(_�5�]�(�5��YX�MAҔ�� J��hı���^�R��>m���/�����1�-s���E�+�S ���Zj��l\<A�2�d綶y-pw�
�UA�4�)�w�"ܕq�7i�����$�ר/D҄�i��Q�|,�#!�ػM�w@�u���Z�xB�"�wy�A�Ms���]L�R�T�������f(O�3|i��E=���lܨt��B�n:2[�U��P�� �D����d����J�ߡ���׈����f�ڷ��mg�Ϲ�r�s�d�-�"2Z�Oض�fKs*�X��y�/�B���\w�WMv	-3�tΈ�-�-<�������2��]���a�/$I+A�~���ה�v��憡lh�.�Iz�x8^H��I̳�\E���4��7�Ϥ��#?� �4³P��~�-�H���~y��6h�G��7%�O/�o�s�*��4�6l��k�� r!�$��]����i"���J#>3����]��l�v�	���F0x��NM[�o�;�8]A?�����yɴ��VsAh��h}�9	�
�'�؈7u������^��k����y���7��7#�H;��%�^H �&	`�W2���	\�c;Sl��������y+���e؜�#a��%�"27CY�ܐn�����J!��U0����Z�\lQ�0�v�2���.� S^���s1����Wx�b��x�����%�*�2�WB-�8~ 7�5�s�Ӱ!L��o�V�	l/��k�$��BA,�K�9��������u�M{o�m����|9��՘S�/�*�At�i�1����H�2�f�T�KAh�@r�f?�<އ^��m�o�A���DL�Z팀tM\L)w�NI���R�,q>\9;���ҁ/����4��ۦ���y��{���ಹY��_�ԣ�u�<$�''��C��O }���b�X�*�΂��*'n�V��W��R�k�7���VW=�)k-�K�����9��4�>�ܦc�j�u �|	(:G�Wń�D�	
�����ު��P����t�ԋXE�ғ��V�r����������.L�\=����ȓ9 eO�J���h��Q��-�r'�@\����A�$���p�mP�������󾕂e�Oe�=21"�S�b�x���Dk^�k\ޯ�[>OxkmKr[.�W��zꗯ:���LuG�gX괃6j���x`� �c�hn�:��su�iko0T�@L94��.���T3�w�M�.<� ���k�q]���4�;��H̑���=1,�`DNA�o�>��pՍM�ĆܕN�J�ƅ�3V��Wo�9���b��հ�˗�����9x���v1�a�B����%�������0e<|4���,���*�靼ʃ�!�\x�~$KueS}�J�(GF�1YP}�AB0�O�T�� �d^򯾬�
x�� ��ݟ������n�9�
)�7
�e�c��Y��Nu��^tL�����^L�f㴹�5��a)�5*��, ��
�S�ş�ߎ��uuv�o;��Z�����P��6 ���:��W�A�~t�$-���K#��@Ϥ��� ؤ(�Hh�1�x:�I�{e�t�DR�;0��lZ�n�Y?��x6E�L��2����Sm\1Lw>\$��9(�¦}����O}�\n��QU
��W�0;J�����g����?ۯ���U�ey��.ج��`���g5	���@vZ�r��P[�obt-�o���9n��DS��=��%R�A��@����}�4.���zRM��a��e^�X�։�M�7 O�p��x��l7r���#����Pz�2���:�k�y�7�emMK�ת�����L��}�]7�>��Ә�ki�Uh�,���1I����L�UIЗn[1���~i>B�`�IM-6;�SYhǯ8�K���%h�ܠ'�*��0�h;]��.u��E���,��D=%Y�Q��[|˅%Ǯ�R�i�H$X��g5Dټ��ˮ�,�t~�dT3��a��w�� �t{�Mǘd�����������J8�t	�h�/i��i��T!�cj�M-o�܋=��:@�(�����a��b������%;e;7 :O,4]�{;%@��z�I�R&Ǐk�c.��_f��r�A����d��?orJF�ʰ�&;�ZG'4���W*A�@� ��$�i�xY)���3�@	�mFp`�WNrC����ފ�R=�Y��4�l�F�d"�21�tYlʸ�"��s� �Ц1j0���D�F~��p�H����Sy2�i�cǞj���6��HKew�u�IM'�~�5f
��3!��Y�j�cX��e�={J�>xUX�;��WG��H���hw}h�ψ���^D�z���W7�`!jY�|ɳ�qp�ao�4\!tV�)������^����Ȝ��/2��{�gM*�t�L&~,�������������1uAS}�'A��$�9�>v��D�;5S��v`��+�roe>5R@����V[�.������0�CP;�@����[�_�+�Ve�C|�jH[&�|:ĵY��4a%Q�d����r�RȼG�2���
g�� �+5��k(�"��F^�H*#ȏ
��@њ�Gʈ��4n���O"گ9s\&�gV��Y�2��������~��Ctw���&�BsZ-jR��{T��@���?QZ�;9Y~�:�G��K�A5?�D��<���ǹ0kM��/�r\�Ei�.B lD��{\���1L�B��e�,(� �O)�7Vb��`�E��R�KN7ځz�7��x���p=D�U�J�z�dx:j�=8O�U�a<�y������^�̛�)q�<���z�y����M�����ԄαV�a;Y���#j=><���`��5<%���379B\�wHF��?��Y�׳�V�r������O�*;�<�h6oi�2ɩ�E˳ �U�����M�:�G�Xi1M�ñ2ņXV,n7�Sֵ?�'w���L��4@�J�oH�I
�>�«�s�'��2�:�.�$�b�j����ݔ]^jA��y/{7��u#������%6?�"����M��UM�O%�ڰ����g��/,*y�h����еBQ~p�i{_A/+�7p{�6�c��B�Bu+�,y��z�j[[(�"��'�p�f�V�9�� ]����te�p��{��R���$u��gPm��b���97�|��*��K���x��V�|&���ܽ���QS�=՝G�����2�'���>��e����\�WB��^����'���)�_4U2���	hޢ_�٭�o��;N�@�=^�+�}I���Z�� ���I��	$)��/zB��﹵���̊y]���#%�Cvn�4 �z�cS�xKF)
h���S�7�bn�mp���j��z���U�H^6��8��М�0/���0;�G�w$���V�`�à�l��_M�9k� �c�*
�]���?]�̔W&���r��~ާo)yd�[b���}H1z�^��5�쪬:R��	���uy��(=O�'�"�lHB��j#	��.P���Ţ6�XDH	J��Ȕ�V͂D�E#\H
b#��뿉S*��շ��r%2�bŧ��U�4���$�м;
H�C�4��h1p��A�Z��"�w9���]_�c�'������2�P�d����|��[w�^KB'>e��5/=���b���+\ߵ��!�D�[�Sr�q����#����EI�4�]
ń�P�'���}�+�w(!�pD��0LP����#b��V��Xlm����!�P���6�ڮuVSм�$s�a_u�X�#f�n��1D���c�N#q���~^�l;󹰲�y�E��1�J*D8�G ������)��`yK~y��&^YuҎ�_E��/
�T^,�,=�&�	�����nͼE�������OUBr����>��~����	x����[�iN��e	c�l�52�j����͙�u��nn��	�7Cy8IFX��P�dв���&���~�А��Jz\��ʔ9�P��]~,�0]���ch���qQ�7\ʛ=�
L?�h�T�5���oJ��h�08����ӯ��Z?�Ñ���6�7���~�,�q�U��NDv�M��e�_�l�.@{mp���=x
�ur��Z�3�d(�/�����7�RH�QA;_�O>��*��t�s�T`մ	�Q�U����R"y^����/��K�-�?[�`t�MM5�]%<74��������'���~B(}�1�沯p�] �Шj������Z����"���5�Z܎�$�]l�&���ϲ��ܫ
V��%}cZ�~f��y?���lG�⋥����$�D�R!,gD��"��:}�$��q;zJ�:�a���@7����\.5���J :�u~�)�����1J9�C�s�C��f�|��v�qT�M K4�8`
UvBT�i����踦�$xܮ��1���@��>�:h'�El��y����}Lz0Dpn5.��̼�aQ�g��������8��Әp�Y���lD�������H�π�MD�`�&��90Q��k�h��	j+Fi
D�~M�[v=2��0s#�w��I߈։%K�+�uR#v���d#�`b��n�V'&�m�c?�a���7�Nn:F]� 4l��p�X�����6gaƞ�JG��-x��=�]u`��8�|�p3%AK������p��mKwo_�E*<�e:𶚟�t�|�X?��,d�,��'V����*�H/��F��Ѻr�WY�y���!%w`�t�\�7z�P�ӝ*��Θ�Fm�#��i8�b��Phϻ�G��f+}@3�L2�.ǡ�H��؂�D[x<�员g�y+�q~d3?�X��}�HЋ%\�]se�9}��U��A�qc�2A�+Wb��Q����(�\�n.\BAgZ���i�Z*	��?ʦ�GՄ ��r{�~w�ct]���-C�����c.Kn��L��K�ȁ_���( �����S�:�Y�D"��Z�TR5#�p���t��wwC<��2�P�xQ|�'��4|mV���vp�v�Ο�I����H���P��mz��x�G�=!~(́���'PC	�&�I������Z/�@x������q��n����up�c��!�Н�y���E��)�X��)J�F� 8��ќ9�+�1˃a�.���m\�:Ֆ�JCE�Ȟ�93�%M-O���_���-Quן��<��?����4�8��q[A�"���}�ϛP0,�Q"\9�@�I�.[��q+��M���w4��4��K��\��G&��K�'��1��)[Md��f[Hk��@�yD���\�����*.�:$���[ٔ��v���h!����j��� d�e�����Ș! yCr�xA�����޾����\+pm�ּ�����:}�],��G`<۞���.���z�C���J�@q<Y��VF'�\��C;�[�����Բ��
Ԃ� k�N�]�J��tO�^[n����,}�۬8�B���o�����=p�A��$�	H�~u�5Fn�]�Z����A��E�Ð�-�o��$�7�ig�j8"L�.��I
�d̴�P�jY����JA�0� ��E��� ꅢ�N�$
J�B���~�@KDx��v��(Ak��[Q���&v��2Ҡ��/bK|Tg ng�+|J,�hn���ku�3 �8^]:���~���޲�wRa8��V>n��jd��2O��{bϕ6&�H��y�jap��G!� �{��A���pJXj�@:Zv��=7(��P4���ؖ��y��bz�y�%���@�r˧a�{3ɘ���
�hV���-�@�����i0�3E�<�k5,����{-(����f�o��*uY�Q�e��h����DIe�]�w��u��m��8��<�o/5v�T|�+��JX3Mq����_h��(a��7G���q�]mI�]���Ǳ�X��e��U��/5�_�,�F{�;<���Jb�:����"�ȭ�X�xb�UV�k���Kk*�4=�
2�d�� �pI���B�20a��kigkd9ӄ�!�t�\���Q��C�᫳�O�&��e�q�8 �����g0�1t:��lO 1znjs����#��F�&
ȏ��`#R���7���ϝ3C���rz偝
)�`P^�{���0,�e4r��p�bf��da�!��h�~K��+�����c�	;>�Εs5,\E݅_(�L�N�� �82e�f�T�>߼�}����;DI@�q$�8E}���*H�'�R��"�ϊ��J�S7в.��満�<���M���S��p��W��Eq!������Xм�3�3�4�@��B��uZF�1��a�����zoi���[�u�h�d\�) �&z����4�ފ���{ �a�[C����(�g��G��ӵ
a���;X@�U5���v088�{V��j�|IvL�I9�љS  ���`�\��z59q�+��0\E��D칸OT�|	��ڷY�H�j!�WM�Փ�ű�Gп�-͖�ԫ.��"FŌs�߈`�M�����!뭢)Kۺk?��,���=����K�}�TMuo�	ɧ0q����c����$PM��Z����	%�����P��G�Ƚ��������3��Tx�5csѯ�d��FS^��.ٙx�Bs�+�V�(v�=N�X��@�z:�/(�<Z꿈߶�˳����g����'�VN��\��ĳz���btאƾDZ�#���^L�C���'�H��z�-��)6�iY�k=��ЧA�fk?w�X�/ڞ ���Q�Q=OKs�.p��-*"�p�B%%�j��<ږ���Y�REJ��g2-��߄y
�w������׍���j.C��"o$�v� ��IP�j7e�_]|�[��ɓJj	k�N��8�$&yA��������Iˠ�r�E2�{�>v�0��P�3SÞ�&�ɑ�������pj_�!�k m����:JHa`�3F~��3�t�Y8]]%�`�ypw��J�$��\G�R����0��xFB�}@��T��0	B��5c�!�"��^'�Ƃú�2�<A��e`&@��9]xۂ����"����.�J ӂm��ˌ�,��G�p��i�CS^�ܯ�+.��*Y(��'q��_�>����Q9�����lz�j�n�	/˺�y&؞��G����K���6��h&Zaa)]d�1	���f�Z8Ӧʸ��[y]��G���ƍW��L�=�9��h}�����6_�����Zǟ!$ѭ2Fu� )�}��zƚ,�Q�P��B/b�gZ�F0D%�J䆗V�qþ��n�Zz�:�g8;�S!q6s�j��heo����<{ْ����0C�"���>�d$}^��띱B���4ű>�3�a�ç��R�����W	�E�I\y2f���F���/�[��PCc#0�ytx�@[I�Zނbpiu@}�)�!������'��X^T?�x�r��?x7ɲ+|���7��e,��B(��Z�]9Y��:'�p�L�׎_�(�/y��n�fѽ?�nr�b^��������`N��i�ۄ��;�ŷ	.���Vb��� �$~ɽWw��h��4���B��u��aC�6��g��WM�����}���u���ΐ ��8m��:��6�N-|�XAc)R䐯���_3��
���~c����;=T����GMx��Kv���3̷̈����ي�ga*"ekj�2C���h�a)L�'{/�-z������3�5�R;����q��Ɨ�����e�"�
ߏ~���!/�q=��w��s��6�`�����j��yD��l��1H�� ����7�Hs��,��eg����׵�l �[Ɗ�5���'��ȝU_����x��ίLQ���_��d#���*&?��#3�9V��D�OFI<�.����g��-Щ��c�X�0�#I��'�����nR�]v�ݕG.�|s��Q���qy�w��bg���C�si�⤐�и쬮��Ґ����[F=7t�v�j�%6�^$e>�@/��38�	7����~)�O﨩N��Q����%�� \Em���	[�P���)H�?ȴ��EG��*�*���~hn����;�
�{��O,C�::�{�mMĤ���V�^����Y�j��O�d��Q���������/��0[#ߛ�7�m�Uv�V���t,5n�5g?�����V�sП�I����J��U���N�ǟ�k2�:�j,�/7ȔL1?)>�))o�#6�@��6So���h|�,K��Ǉ�e���<�	������˷n\��Y�,;{0R�3dWhn��h�����ӂ�������d)V�Ut٧���4��R�������v�U���-ïI�M��
x���؏��*v��vK��#���q{nL�b)��8�lO�}%�������O#1X+H����E��Q*�';v�EF�,:D����O'l L_�Ҧ�V�W����m��D�矻1�K�_}����O��v��L`�}��r��J�7Z���A
}�Ic��eM��i���Q���4��'�ݹp��D���"���=���W�&���~�tX{7��KkԮ܋t��i^�l!��)�,hS	��X�l�+�����i���0"�Oa�$brcC������17�]H�n���B���3�c�0�����G�7�V�s_Z��c�(
�<�?�=��~����
ըR��<�Pq�ʾ�8����w�#� ��s|t֫����]J��Q���h
Z���eC�I����#Xh>�����EҶ�lH�%-��Uvʲ/�j�+x���K)��4�,�Ka�����L�%s]R�����D��HK��c��}�Y�.h�YC�y&����.�9����zy����VrI��wk1��0ɱ�����x_�S�zƢ�ϢR�'�DAH�&��<�w�`J'W�r��tM�T���4my���K�E�M��D�\?$	NM�ד�g��NrGM
�V��
��o+���@�>�,eB;D�ށ=D�7е�r�W%P��&\�C���J+ H9�:�`Q�p�]s��9��D��)�����KW}s���e<.�}".����&Z�+��.�᫞���c=�U��V �6�@?��LF���ۨ{��@-Dh`���)��_�J�	�⳴��_�K��z
�xn���'^G�U�#��g����I_pg�\y6$�	��_Q�vWf"�1H�j&[�>/u���R
���(p|���T�yOru��xc~2I}�3�-����nd3
!3�yN��7.�{M��ɯ��x�מ�b�2h[.�1�6�������_XN{p�j{PHCWZ�ʡ�w2��,(�A������%7�b������D�JpW�*�n�Rb�����a�l���	ڛK�v� ͱ2��y+V_f�~��E�L�O���-I���GK�ˮ3�*��.�Ϊ1{�׆J����"��+�))D��~\�2��g���6�T�>�b��@�M9c�:��/Ŵ��x��kq%�{E��@d�&����������=�Ь��̀�5��t;&j�sw�fZ	Lxr�������:�1����CZ�mr!>*��l�LU�uo��b�:b�� �)�F��!
�8����P����ƎO$a1��$�˷$ru^�=c� ̘�;�n�N�ǃ�M�`�r�9�HVm�y,,rc�0����3�_'���-��p�MɄi����q���~x_&&�����Ki�di��t�9(	`A����rH>�U��c�Op��W�G����?(��D����p����Q��#l@ö^^�����ҺK���k��A�+
�X.��������f��L������i��юp&�{._����m`��+�1��-�w�9ϒ�} 8�~��S��d3�&��(_\nkpi��8b���밳U�u�ݗM�͒}dK��G��	�P�d���q����9N�F�����tA�9Mr�����S�$��^����� *+M�T�&�7�5#�G���p��1t3�Q�" c���|������}��u��A� ᣸?��8O�'{��,���9&k�Д�����bdh4��+�tSmMے�����8J��N��0<����K�����.�9.O���i_�ٻ| �̯Z���kXw�
H��L�,]d�ps}��?��`!ͯOf���(�ʒ�p��`R��h�7[�>,�S5����s�J~���������ƣr/���@`~�w�Q�kX��sJc@쫬��g2v��Ϫ�O����Q���x�;I���BFX�jgACeS8vp��"[N�%o9)��"���c�vk��I����k��+^�p<%\թޠ2�hR�=-W��m������G#���u�"��
�+SɝOG�v�H�=T�|��w�����������3�6Y�G8+DO�ʄ񪌥�z�k+�)�ר� B�̷����| �o�9�rcк��D
;�w��s�~�s�ZG;&0q	Ѧ��Y��Q�|6�GG�Pew`��HIK���p�:�ڈ� �1􏡇Q��v������ڠj��~����S·qxb��_��F��x�;~J)&���˾�U3;bc�=:��~��G	��A�㼥�Aa���ֱ�UóU{fN�����j
���c/ԇ����9�b�� �\���A����zƋvj��eF��*c��x� ��aXj�F�~~VQ�)&W�|��Ad�&Bay�)euwN�������� ��j<��Χ%i��`����p����1]�?��5���pw�w�5���~��,s.�6WIO�3�J`���mA=&�l���US'L�<� ^`���q��?����Ӊ*+}2,���0~V�%�hs:�w�ϳ� ^G��~qpb��	�6����(��mE��׃����V��`�|9�r�icEk"�H�⠑�T�UZ#�F��
��t5�qW�(ZS�Z���"�b����J�g'�b�9���W/CL���<;�%[>��<t�gOQ->;6�\�@�!:a��l�/T�Tե�IF����0u�:^�'$�P������y���w�8l;�k@���İ9^�N���/��'N�b�����h��~��6a�s�h��Y�A�埭�6����,5�%�b$���*+�#\|G�!#��xS��O��3��)=�Й�lQ��CI<)Ӣ̂�����rD�E��8�s���	��ڡ�aHM�Q�r�l.L�i���Ec������7��N8�	c�T� td�����v�<�"�az���<�ɺȯsԕ*4Ƕ�3�$e��GO݄c$�nJlƳ +�	4��՜ ����!�dN �G�[� ,=��߽�Zqa�I1JQx�|�%�Jz6#� L��o��K+$8��5pQp�P�"����ء��?���"=!�R�	�L*�%@`�t��_��?�� �r���"�Xac����TD����+YY/��(���#�����ѐ�O�PB���a\��Uƿ买�+W��Up�#��4�|��dy8���qڥ��)��a�0�*�!�ڨx@�o����-@N&*10� ��Ub�S��ZG�}:�dw�#��\��s�GN]�G�7����.����7%��D'@��:"<]��%��3k@���N��vrF��a�G'5�X��Z�vVCMԖ"�y�6<*����Sxb_6�|��y��4k}�{�ۍ:P�QW�v��̝
N��9���*��tn�^���2D��vDķ�`5�r�_��'bg�ㆾq�4U :"�� �n8��ɡ��]��9��QJ���(~��e�0��c���'B��ʖ%�^�\��?�����\�N��f;+�`q���,��@ഖ��X�m���d�����W,I�U�N�@��Aq�K١�����J5 ��Xk3��t�������0���s��j��N��+�
�4t��\�����)��>7$�`�:�=������y�P"�����PU��k��?��*Ĝ��w[`�<un�����:4^��չ&q��
Wz�����[y)�����e�O���������?�=����olʱ�j�t]�:W���{]ٔ�Й�����h�h����R��n����.���5,&CX<�g���J��da��:��;xe�\R��c ��m�f^$}�G/�IR��4y����0`��[�Xz�d:��D
�nN�D7�.Ʀ���b��ظ}i9O��O�Й�O�����*C.��.]w��-ɤ?���E����7㩏n����	����tv]�ޝb�	L���	B��LWeYj�Q]iQ|��ˌoC\�4���\��d����ז��ty4�~��0rΣD���Et@���RG䏥jf�ο��CR�	�z�2�eĸ��������Sq|Y
�g�	Q�'�;e��'�*��&�M�q`}Ǳ���6���K;���"���1���$RwtO1��o�X���_Ȼϗ��O�%�(�6������-�b�QZbFs?�(tC���sG�D�s=���R�l���2�'۽�	ba�=Vdp�n�En�˦ߧ�HǤ���Y�w��}�bM��`q�����U��U�}��]�4�1�
<��:��j�T��(ĀER:��e_�/>�j�=�[�d������Ǖ�l��J!�a@��w2��K��B�,zQ
P���F�3M�Y�	���;jكt
:�^|!a�X���CA�!�!� ���ԃ]=�>g�J
f�۞�'͐b���2ɧ��%_D������a�>BƁĆa�+w����W�H�x!�rem=�R�&Q�⛼��}���c�5W���+Xu;<]ҴI�*6�M9�j�7"|��D�f~zT4i݀��y��A0�������c����8riէ�:�ҝ+JQ	�� X��ɲq)6ѸSh��O{��~�E��y�6�KDh���p��������s���J������#� _��):$�#��y��>x�^�}�+K�OD��M��a�RwM�T�̅5c����S� r�M���c��x�Ǒ�:Ox����m���Y���w�i �Ɋ<�@�p�w���ɹvD��#�C�H�0Q�xJ69���Ip�!��D���z�oq�Mi��rD�^��'o:�._��k�;���@ƙ�k5:C���j�Gf�kYm���g������Rm������� �0 �(v/����Y&����K?<�ޚ}�?-�y� X����sO�Ѽ2������81+ۦg��큀����uQ}����0d�:�%��E(����Pq���X��b1���I���P�@�۲��=E0���aʿV
۰���ў`�!?�H�j�RAd�0���9��� �B6~��*�Ws\����W�z���^�;��W�Rt�༒5�V.W}uK^o���dy�-�MD63y�j�@��9F��k�Ha!�yw�m���0;Aa��hv�y �UC&�h /����߫�H��,�8p���&�y�G1)�]ۇ�M�-H?��Gpv��f�#���L��Rh�'Y֔��XU):c�d�wN�r�-պ ���+����$�P+���N�of�&��s��~�P�7���VͣA���72_qg͓��F�u˩4-Y#
���K�{C�mv�ڊ$���P]�]+����Q\;Z2=r1Iolp����c��?:�3)8?�C-�^�_8��g3 �> 6dOk`��
����3VFҿ~@�g�#��,��4���<�ZL8[5��6�P�me�qg'a����)�7�>�=�)B,Ŝh�ix��O&w9��Ў3�����U�x�8^�|@�O~��ə�������������#�p6�c����65H�5����^��d��ڻ���������6�/v��I��-�rK}�0Ϊ@^����\����!�E^�x��1ث�t�s�j%��1�Ad��ǥ�[�N���]M,=!��Ԑ��(�ho���l;-ATr�3^�b�.��p�7XZX9�+ߑ���ܱL�N^���t�p�TC~�[�2]
�&� �;�ك�Mx�X���{��i!U=��'�2���{A�d�L&U�_k��t�t��W�t|���r�V�}����M�OF��) ��qN�*��ω�ab�[{���M�1y[q_J��Gf/�PAٯd����������"�z�(�D����LR��iZ1���e���Xk�v���;�Q2�ح�v�"��:��a���:��s1:Y�õ�"]��2���1�tZܚZ'�=�h�r�ު�)�t��Jݭ�W���/�x�����!�'��-�]�b�I�M4��3ƹ�tqOQ֒~��&�= Q�I�r�T�̭��ˌd�W�O��q�H�B�uS�����[�����IzK�_�|l�R�-P5�t�@����#��?��|����ME���q��kP.�$���,�CP.+X7��Ye��eGә"i���/Z��*���������ѝKČv�a��l�U}�_�#Q� A�q0�]���������A'�B� ���Qg�w����+�SN�-�a�b���k$GM�D�Ha����^���� +��tˆ��A�����[Y���r����<Ui柽yH���~@�����;�T���րv��L�O���gEu#��:���@3Pg��ם���	
���Ů���.��I�*qD�%K m���ͣ%ْOO�mw�6�J?x�e��Mxd@�ؠ��)~<*��رp�J#9� ���:2�8,$�é0s���9�6�k�$4?/ݒN0E�t壺U��h��!���Mo��	vǵ��,Yn���S�h��7��|6�6;S�_����G��8r͎-P(\�����@ǁ#3�Z�x'w��BM��PfOb�/>���)���e���I�y��}s�:��'K�/{�Q޴H��ϴ�Qo�~ 9�9@�ΟhZo}�p1�>�Y�Ɂ֓�mV���
��L�:�,w�~�(-�<l��}/�u��x��F����%�o:�����I��>w���<lk`�hS�������2��Ғ�q�+r�RU�?��Z���%d*M����Y��8U��2�K�%�B��G�=�������a�gw}��\Ϯ�W	Q��&�+�پ-_�}$�@�#%�N"�<FǛ�g�n.?�o{������.�y�:-/��#m���Uޞ��'9���^��㦴�H�
��߸�A���'j�y��$C/3�WN,��|���R�;�I�<M�B�����ט���xI3��Z) ���O���Za��(�d����$�4�`T�L�OU��"6�≣�I,��Dn(�=������w�p���D�Q���2��G�U��ܙB#�oG66��t�%G�l�XA؆�����o֦��8z�J��B�$��znYwHs3�Yzqw�#�� ��g����B�^��q���*�^�/�q��c�	�A$�a�j��{��u>BĿ}�Z��2�%9E�XzR���y����,��ͦ 缜��Hs�҅��\��.�CKmS#�j���bRs��F�fI�����Ɲ��'
�&�Z�����C���?���NrX�H���Άͻ�[���ZO���@�H,���	� 8����_�PhF�U��\�Utd�� ��`G�
����ڟv�l;���-6�㛚Z䉱�$s�Ò����o��_`�t6T)��i}l�(�sm��@/�+ug��(�繗�m����*E#UZ~�h, ����޸(��-�oe2�%�p��.E��vOF��w�%Y��k����4�{JbɃ?L�A7���o�v��f�L��"I�9����2P�V����:1�=ڿ�YΡ� �nƷ0s����x�^i�����6=�u%#�l��o<b�!�Ṙ�¿t9R�0�������T��ɒfO�:�Iwȹ}aF�ҽI$?�g����<�]�:h���QzaAƈ���#JT�C��QkX�3�]������z�����b��>=�9���w���q8�2�3�T��u��SGs�G��.+�o�*�#����62(R��P+r@w+��Ψ�~s	\�EzE�<��?��&���ͣQ��
�O� �~f�X0�<ࡉ�����A�Vc'?�CU��:o����n���M�����)H��hI���'p۽ϭ��Q�~�$hoB�n��p�@/��(���ʳB��;��s��K���3X$I"�!�'-�_u��{�3�۰������N��h�����>���'��u�t7���2��Q~!$� �S®��#&_����D�}M�0�����S���Ή껑3��3˗�ϴ�`���f��P2���HR�'���������/P��k_�Y}V���NT&��NYpb�E5�M�E�� �d ��ʬ��y�,.TQx��6�'�:��:�e`�6�,E.;v|Z<�Xu�����L!>�K#��f��ZfA5�3�"������{�S���c{�(��S�����֥JHT
Ké�(��_��������,	?�K��L��]���_��h�ě_�2UY>�	������ʜ�����]j2]��P�ٟJ�d��BS������E��X�P�ܮ^ss�@�1M1U�j��wo������W��d��C/ӒK݌툗���ߎmTǼW?�G�ꛩňG_-���N����
�2��e�[LP�~7SU�C�J��]�T�R���"3X/�7G��ۮͤ4�?vm�������q��4崥&}����6��z7��GE�"R�4j}�@-s62�Y�\�$����I�;$~�7����n�dI�m��k�L9b1���� ts̴�6>IJ�:��k����<3�ޡ
0�S��O���r��ij0�*�:	��R�oi��F���؅���Q�̋	����X�
�űڹ��1�y�n��A�'{�:�I�4��a6�wI�>F�c�N��~�O�f��~��~ff-�]q9�؋�<o>��U�k�P'�Fe_k�H� �h�ӫ�t"}��3fE&���1ד�k�	��pm�W��K� Q���=H.RS ��OpS�Բ%��D�r��X�����ߛM�)Z�O������BF�nO�ў���?�^V���!����߲K��ͺ�hQ�gJQS��E�������qepZ�l9�@qq�����_�g6���ժ�K�yC���r���_�+�9���7Tۅ��Ȥ��w��1߃�&m��1�L��C9!�-��| ��N�]R|���v��`GdQ�6 �Ũ��	e��$���ˇ��ܙ�9VS�P�Y̑��U��"c=&�pQ|V{/F�+J��o�@���!:b`��IV�*Ĉ�ԂZ��'�؆w傱j��{\�rM�K؜P���# �D�U�4�/ehk��)[�z�,�qx������lN4N�ٯV��5'�D�S���{��2�NF�@��YR�?-K�c�#�a��t��P����o�]v�7���
���nk�0���!ә��T���MuyL#�k�sOz��`gf��,�E����U���D��ωy3/,k&����U�F�|_�X����}��D�L�%#=�e��SK%���oRK�^����Y���o�3l��''g����k��N)�)�����}�l�bFfYd5U{޹��Ys�h�zڗ ��7`�ǿ�'-I���PG�I�M��s4�c3��$1?I�(���"|3J��e�)�"Vh��0õe�6���v$}'�����	�3h S�C��]U��@����6��Nws*�S?��h������1���KJ�-x�����Vz�P嬚�����o��/&��e�Aq,Z�E��q�	f���>h�;���.!�C��E^ʉ�b7�֛'O�Ѝ�g!��j5|_��n�̜*uk�K�	����h	(�&�q����`<��w�@��7s��d㣾A_�Q����K�Cz��<�/�cBxm��7*M�ouY<�O�e?�=�=gV~"������'��� V1e�F,p��!����P��x��0�ƀ�%)�}�*�5Rӊ^���Qa��{81}�������OZ����j��"�)��&��hL�	#�E�Hd�T���o�e]/_��:�rf
5
�#���^N`��%B�R$�6n#b>Ƒ�GgU�2uR?�|q{�����m���Ng,�a Z�8��z������\�3���'i�R��p�6�^������y��w��|"��l�y��껖E7����b�����b�W���Ӿ6P�:�6�f#Œ��\��L8~�S�a���p�gū�5y)��;� �Y-4��ٴ��˹n�7�Z�eJ�9k����x�mlF�x�J����LD Dڿ�J���G	����D��<�V��Z|�F��E'��"Q�xb�#k��bd̃5]hcK�@�(�U��3J4�>�X�j���_a�a�����W��5�)�'��*��S(�����D���F�����Bz����4�݁p�G>�I܀D�eW:���傑 \�΢\���E�-ĳ9ؕ�aM�����+�	u�J�wde{���������8�֩~��8�[�6~7Ņ�f�V������������1q��3�i�㹖�2�8R��R�(	���Fp�tuB�����z���x��,N��>����e���,	o$���ʲ*�Rh��4SŔ6�/C�����ʹ&L�G
p��U��Y�����fD��G5w����r�8�G&�ft�a|����j��<(�L_�Pր��W��_٬��l%�X�W�-"|m��ށ!�Su0�}���e�r�O����/�,0�4���u���?�(��#��C�s	�AN��/π���~6ށǒ�=Z�8�Nz"'h���-7D��Q�"Z��[�Li���kz��(&�ѳ��׺`_a�VZ�;R&-$eD��1a튥��fBND�_*��������4I�'��M�����W��U���3����h���Y���s��] g��:)W�?�]̗�1�>x� �oˠ�F6^��hκt+�S��j�9hr��Ѫ�����K���]H�^�H�v� Գ<k�U:Gx�9P���Ɖz��X�t�����*8�@���9n�Ƨ<�($��d��Hi,�-��W��U /���k�Eľ@���r@�l�gVLmgJ{">ì���d��@��/�Z�f�Gba(7�[��YfY&�^��_�ųU��ށ&yR�<]��$2��ͣ�|�m��>�A.��6B�ܯ�8��~Mdg����q|S�Qd2KX�Ѕ�&��iDɾ�C��6��m�TƉ��Q&��ͬ�xlh��\��M/�{Yrw9|��b����v���I��iv�s�ܶ���W����դ���j\Q?��,�;3���ԸA�x���(�eD.��캿�hC�ab�>NĮ��%���7�CVi��g¯FG��=�<էf�L�wN_�Mp*��ʥ9������[��]q��5
�~��y5�O 6J��ZQ�\DO �q�����]Q�	��)Y<�鉺U�5d����8��Bn浍=��!+����:��9�-sPۻ۝�cu�KO�Pc��ҡÌw���kXgB�!�0<A�?��I�P@�7���";QrY[A����'��߷���C�n���_}�܌���&Ђ���~�Nr���ݮ� ��l�g��Cg�Ȍ���ZQƳЬ9�}k0�g�c��	���59�}�5�KV�"� ��.�82�FD~kɊ}ʦ���ߧ(��77��6�U1���k ���k�
H�Uy}��B䊑�t����� ����/��cXph5 �(m�yE�p^IT��8�g�
)bg�CՅU0�N���l���%(ND_ ������6�9K��F}Y� 8��U�NNd">_#�3-�A��f|�$�WP�!�݅��+��1�WȚU**�6�v�K��H���Z��lb�.ʫ���P6�T[��fuƕ<�=X�;h�s��g:���V��7�\E���d���~�x�Q�����r~"l"}�}x]CQ[|z<����MX��T~c_&�e���E%(��ۥnwr6��o�z���+.�%�b��b	s�*�w�AB�3�!�:tv�w�j���b\{[g6&:�r�M��,��Pz�����	�!m���2�^��*�%C�6Td�wS�ÎhZ6�G�އ:�p���>X{O�ajZ�aԏK��C&��<ImS诣n���r�$g9�,�}��LR���ߜ�d�{	���AUjQ�4��P�-%��-����>�}Zs�'3 �ۥ��W#y=L�X����ۂ�s�J�k�y,vH�1�
�7}Ac�%����K0��.t���q�Cat{V_���,��F��`!G�g���%���ZF������ Qء�p6ް��+b�����P"k߼��e���7���F�c���&�T�.�g��da�U���RhY��ƍ�ʹ��1�۰h����J��R�ù "�E[T~l��3kb����aN��ש@���
��E<dYʊr��Τn��>LK���<���r���5m�N@4���ьz���S�s�r��޹�	2F�1��;$M�;h����g��/wLR�,����Ɵ�t��ksE.���{�,�ˉ�gDC�r���ɥ�J�7��b�(��h�lA����TZ �	��V9��Q�p�
�{ӂZW,��;�Z8�
��0�;�"�
�d�F��'�����9����l���q��HRKI��l\,阯O�<�I�zkJ閸��V�*�su�eǠ��3[:RZ�E��U�{�2-�lb`����F��O�j�J1!�g�d"_��W�.p�,m�}�}oA���M:��I������GR&B�©2��+O M���ɽY���1y��]'�7�w���'⺚偷HJW�u$~���כ5:l	G��g;@��u�H�yz�)(9�vl�>6�Ĥ���W/�ڑ��FQ��a�+��v�W���.��y,�˔�W������}��r��8&N�W�U�:X?��<�@�$�K�����Ԡ;?�$�^-��/���r_�2�H���^%?�(�J����:�	;DT^RHۙ��ͺ�qٔn�ZƇJL8j����צ���\����I*MU�; �w��@�M�CsW��d�,���;�yWҔ����2�����z��;��5^QaV���
����r�>l�h�q�γ��kP�nה��HZʏ���]z�ɉ^�>�yB�+/n��~��|�&D=>~�	����}r�f�P�Cق"���rA]����I?��(�<8QU;���α��-�s��FE���k��n����<�	�g�R��>��?�r|�uȘ��@�E�/+�i��[t�V�ˆ�����ޝ��8uZ�5Ħ�߭��FkNL�N����?�2'*tk��51g�)�i]��x�G{}Z-���:��f����� �Fw��_������y��J���H��C��Z��:flk�:5���:CL�
M�Jf~��h#ϸ��L,�H�|a)͙2�d-R��c$Tb��Y����g��ߣ?>���s@<z4��װLEf�d�E��1kS��Yհ�JmY��
)�o���:��	 F�v��
��6Z]��?9��T^6>pߨJ$�u�]w0nb���w��3��~�|��g�7���&��Ƙc����L��[!IsA"�,a�Y�[ 0�c��w�T���C�?���K=�ѐ��Y���)q�I�i���:W���z���w�^�hG���p�]N~еc�+����Uw�(�ˑ7�lژ�������"ul�(U3�Y]@��	���~CCq��;��1���@K�_dV��A�`J#���:fw��1��d#=�����ׂ�v~�H�ƴ�m؎�������N����d,{��,��Up9a�<=�1��Do>��Τ�qg&e���|d�����puw{ʳ��Y�#����p\_YYJLϕ�a��dI��V�gP�a�sy��|�3.V!T�osk���HYǨ�cf+�6��0�3��Rs �M�A�M��4=̗�U*V�,��ɺ��]��"C��e4�S��iiF@��g*\:�T�ǥN�hS���u(4$Mx�y�|h,O����¸��&ڣ�Z;��}-s����f4o�

�W�S����B!��I�������A��h+p�$�Qn]����ٖz�[�� {-F4�Hh��%#��'s�Q���?=}�.(ٵu�8(���O�ښD�����m9=��G>��]�����qhy������S5t�V,:F������dA"�YG���?
��q�]O�z��7wu,?��_�d��	]�?P��%M��
ɭ1:�P=����*��)����@I�S(��1A�bV)����K�^-W��;���CqH���H��������jXs[K�*5�\?��"
0٫���7����Ƌ���X���{{�Ӥ�Gȭ�e�v�7]B+ ��ڼi�_P��o��[2�VnY�S��%��ԍ
IhlJ�nc�e�˖����xK(�����1��lœ�}\����aO��F�Rk��P;6F-�I�WzI�߳ߵ:�`yAYP�z��92\��4��p�l�g燕�s�g���
��5��	2�C����\�^_Ğ��Z��@g���ˀfn�!ի�J������\�f�ԟm6*���==Z��F���z���ˋ9��B�]�?�_Y�@�>�A�Z����~m��ԋ��~m`G&����ռȰ)t o2c���f��{��YM�>SP�Ur��hb>��OBN�z�h�������7���CT��Ї�*{�#H��yx?4W=�a'�DBv)e| ���h��kR�;L�ayڼ(����g��E���`�m�'�� rR�㭷��]B���sr�������bs�r����q����I�Q8r��͜y4]��{�L��zr�ڃݧ]�E��[��u��q+p@�E��y���q�{7{(����1�F	YI� �z�wfB{3_ч'|l��$����eԒ�)�sG�:;3(ӈr:ÿө׳wFo_��O�&v.�u���S��5H������G���)g�GdCT$����#(G?�x�>?���+^{���u���Y'5Xk��N\Գ8/FD��Cf'��4�o�M�O�鍑�[��ta>��y��ҵ,ӯhY��c�ض�de����^��w@#Fɝs��8Q��q=�I����J�9o�*������AT���=��|�/lge�vXaZ�tD=�����m�*x�+Č�����T!%�o������^�P}]���#N �z�)��6��Bo�U>��<@,�!���L��k��i�qF�A]N�Or@�S�[���xJd.�d6T#\�C-8����r�#4�ϹNWm1 ��sE�����0k���.d�'��MZ�/�l�m�J��,�i\!�r]fpC<� �ֽ��Yҋ8S�� @�����B��+�����U�}	m+�3�Ļ�.�XQ$ܦ��F�w���m��M�r$�Q��[�.�;t]��3��sy������e���S���:�5f�kh�0%a�uH+C��^{Swl9�NԦ�xu���{�[dХF�F�C3�I�*<6�h��;�}N	�4���AU�SCJ�ŝ�V����s'����?P6�c��� 70����7�l_��CS��NS�g{�5#�+
G���E|�<}�wQ��y*Q�?
����i�yF8�F'Yb��6
���a�}�H�� L��"��ekA�v3�۸v�צ���RA�vK����&��T��@���۽	��r"�X�n��Ȥ��a����8�S.2Хv>�F���L�aƢ���[���{���r�?�bZB�<
�R��EE�.�P�!�qwF�w�*bs�.i��tf�������:�:>ACH~�}�d.#)<�hF���x%MwL�T7}�x�%�"'TYb/�)�$��2IҢ��m~����W��D�>�M�̋���;%��܈m~=Y�dmw5��`;J���d5�s�楄 /��7!��[���Bb�0(��Ee�4
=��I��U�^��)�>}���O1�0�Y�Ǫ\��5� ��D�#������\KpCB���=�/�%)�3�E(�r��R�!M��+)(i����-Ӥ#�qw3`���h�%ig�e������>��g+)���9�����̢�Q� ���|籜����Q��ܨ,p�X���m��3� �Hvѹ���8t��J���Ǖ�ӿ�q�KL2E��^�V��
�Z�^�ffã��y�z_��l˲��Q���#i.�~��Pm���ս���{6�px �K�瑥������ "���o�.��Z{��2z��Q*�P���Dj���'S����hJ��<�A�A�� *9�_��V�]#P}n���fOx��ـ���x?�x���S=f����e��M]At|�?˦=]���u�J����M0h��E�t
�&�d�S���
���q�l�l��׮W�D�#>�#x~]�Z.������U�4�,��*;����׽v��2��
 1�;�;�����)4��nۦ@'aH�����+�KDn��;�u�
�:�M,���c��oJ�&�I؎���7�9�@C��X�u�n8�8a�)�%׽W����Â�Y��BT��eа
�9:���t�(3l�m��j�R�N&p3��~@׋guB��m����r��¼r���~ʒN���2V��W�z��9�N��9� �i�r��㛖e�'��e�Qq',�y�ݪޅqpo�ZI4^��`��V��~��Y�`��ć��,)�_fV�y�خ:J/�sӦw��&zT����,\�)�T}��F�r:w;G�v_Fc�0e��<ӱ��?�T�,Q�m��1�a���,o $�������I��^�x�p������a�E� B0�U�|��Ѫ���c��6��/Ü�ε�U�1�l_p��o)h���N�a�a� �A�=���6��7���S���F�/4��lqI���F%0	��$W�������������b���I�O�����N��`K�Ş�\-��?�M2�/љ>͛�Z^P{�����޴�?�ee�'�z�@��PYPE���i+�������k���Y�c}l`��,n,�$`_�D��c��La_$Z/�˘`�ڛ�KL�ɢJ���))db� Vm���ӑVr�nDAU?���D�]]�yap�ʯ�*� ?7L��+i��T(����)���jע�l<c�$��<^ɯ��M�>�1R�4�4l�E]p����Z��u�k��`86����:"�Ro�==-J���%겷�^�D3��_IvoT�%��� %t�ߊ��@-��6��/B��W,�KIa��f��@��ڴȄ�;	]!
_���^���A��x�BP �?v�m��U!���B�@���#lͶ?�MFg/�_H��tGVmzO9��������v��]�'|L�,$2�0��S���{"�󓪯[�V[u<��񥔊�īrRKz+&�����wf����zș컬�^��<p����/�ִ�WТ���#UO5�Ưc��ۓ���Vq�Ѫ�!��͔�R�5��K�=��aZ�v�تp7���A�$wh|vq��Z��?n¸��k�a1ժ�S�<��k3�4�
7dΠԢ�����������Lw��̂ھG37N��ۡ�?+R*���,񅼾�j3MKb�O:fG�c]q�����}2����~>f� ��` z
*�?m蚬�R�#��#�C�����"BJ�!���'�]�>1��r���3��a?�608'�#[�z��� �ݵ5TE����l�2�h��ύ�*���,��+��ZQ2DO��=+�Nɏ��e�`PU����$`REjj�8guj��?��˹$�A��O=���HƮ��~�v%]J-u>Ɯ;�x� �Ͷ(��R���q��8�AE�h��tB��+Ԙ`���8���'Q[��\|JIt�ғ-,����|��?g�������3�����g6 T׸ U9��S���ࠝ䱂m���C]�I� X}��ͥ�����:���?����O,�~��G5d��oF�OC�]w����i�\:g�L��2?Fe�v�|5�����ٟ�	sS��ş�����.j��ҐG#���,΋d%�~[O�,�B����#x\��Nyܭ%��5��6��xȀ^��HeJ;[�¤�G.ۗ�A���w��c���q-.��\�Ȟ]�ʡu�P�I��D��Ad�kT�3�ʷy\6�A��K/�я��&z/�!'`c��@��;s&8���I��w��l��c�$�̟�lT�Q6z��`�V���!�غ���
h�V����m^M9�6�������i�7��7�w��'�s�#ed#��E�,�ő�%7?�-F�-�$d �|w��x�)}�,r�BnsLВb���?����h�y�f32nF%:H=�C��%��)3��&�ȗ���&@�h>�7��k2�D{���l9�����$��ܳ�	�V�����-�ѳ����LТ&dʒ��R�bo��[������cLq�.�ak����0��v����^�']gw%	˕�Aj��@V���t}�V��
k=���U{� �����.=��i)��i�m��)dWvh�)�s\��s����ί	9��)�*"\~������L��o?\nL��}U��'��mLt���I��CYc��`�ɃA��<�\�yEj���˲7�mzH�Π��H��2��z����x�Fl���dص~{��#��SI� ���h�ŀ�0�$��5�ſ�qzK��*k�}��jCA�����sW�8���eV3��el2����Z3F�k��m������߿���~ԈU[�|����X�>V]� ����B+;���`%���Y�iw|�� ��Z�3�U�7��չ�
~��W���{�[�B���Q�;�ޭ�1!�&+(���".�i̥��`�]1�@�� �5�i�96_,��ტ�f�/]f�'ok�y�w���[U��ZO�Ӆ��tl�:vU!��;��t�n-8#ۂ(x��L�������q�Qt��������ho`!������Ð�E���y�6c�|68�$�G+L�Sx��D.&:z��ߘ�*I�!��phf����gѰ�#��FL7�S�+�Ir�omAª��V�D��*H=z.���l�y�~��K��o�V�aW)���ĩ��l<�a� �?�vG���)�K��Kuh����s����x�t�ŋ4I��$��m�ө����Dp���k��bU	�R󻯩73q����+���b�����Dl�:8ʭj1?��,�3��=]d`ʥ_i�� P���|�u��G�VF���ւ�z8�����_�G�` {� �~�����,FT�*����R�@��v�=�%<���TN�'����>����N��:��(OT��P�����x��b���Ka`���jrG�!)'mƳ7�<{��g�3��y�u��WH���l]�%���ʣ�Y74/|)SA6��0�	尽D���g8օ�9I�KV��Gy�����^@|�_�J=mj]�.�gcUQY5X�#�[ u�ҝ�AFC�>��餚k^4ء:���R�����)�Iy�>G���+�Ol1B�6ݷ	�����'���v]���L�	�$<���a�zz?]&�ob��=� ���`� O�'ϙ͉�����K4g.'�-G5����q#-|�|
l��ujE���';��T��k�KV��Bv�`����Ow�&���&��PVzP��]������e�s��U�iB��4�k��g��J�������0YR3Zj4��|%ńٲ�[ ml�N�B��7zp\+��G��4�I����C���8�yRQ#n��k4�����^����Og�S~v)��S�r�;����e8����Z�٫�Lx#��)R1�ò�켨37N6�"T\\u��V��n|BZ3To6^�+�P�?H��^�� �\�9֋�&��7��A��`Z���<���L�d�b��˙�X"�]������'	��3~殔�,�V����I�V>/*j�?7h�ދ��{��(ٲ����(,=���);@ESs@ĸa�%d"�X��LwoFʶ��s�Q~l�⍽h��
��EJŹ��T?w!|�ĞėN#Q� A�����w�ҍ�cn	;���4f���<�P52���8����A��o�����h�Fi}����{�v�a�[0�ώ�Gqq_��^�}��$��㔖G2'���H!��m���~����o�Qr��rf+�v��[�/˖3�{(���^�AO_9������h;�_�&����]�p��v�����!����Qo|�HOUna��}%��S/��j]be��b�+� �aYZ��䤑�T<�>�Y.��l���k^�zh�Uwg�t�3����X��(�}2a�Ҕ�Z��fg�B�b�T���.��F �C��iП��Yq�U�8��Xs���i��D2�UӴ-
t��q��)����I;��@�\�2o����W�m�����YG��ľ�o�K�kb!%\�p��j`\�<�d��r+6H�q���ت��	ӱ&�f+�҂�;m$ h]Y���V���@�*���2;/��=x�[�6�}����I��Ө�ܸ��f���E����͝)]G{	� �2���hQ�� ���Vk�X�r�~hk��\���-�(=���EO�Z@�]�z��GsǏ1e�[J���R���mz���ׁ#Z;a��e�5?|��$%^;Tu����Z�^
_h��x����(g[�P\��4E
$���Sdク�8�l�*A�
r�7�
�\6�9|L�œ�$�������^�yѳ��줅�����8��ﵿ�.h\�/��㪱�vM�504! �w*U=�V��R�IO7l��/ƀ>L���lW�\�(�� �v�c�]�4�����&r�y&�~�+�����Y#�|�I����UDE�П>ϋ�x��a�a L��5���}K���8�٭��GU�'��Ֆ0>�4�pg��/�K[�r���o� �?1_������M��Ţ�`.Ez����`e��qo	X���ǻ	��QZ�f~��M�x�\�j^݃sX����F�S�/����aB|�I���\��|�_l��aI�/T%e9�-au� �޶�\���Y$�>�5������Z��!�KGY�͑s�l�Fd�`���Fr�8?��a�o�'�������V�7�tR�[L�gu��")	��G��FG;�cm+ �K!ßI���"�t�g�������RSUі�"��?���l�4t2�ه�q�����wߝ'U�(�(�㢰71=n˴Z�S��A����Y'(��dk`�&��o@D����O��P��v ���(����� E�:����,���uyʓ���AM��o����_T�A������-k�F.�\�7Y�7�˘���1�8F����:�(^uov�ر�΁ܕ#��UdBA6svC��94�<�=�u����ܦbм�������p\�B��aS�f��ya��у��^�D�;�nJ:�4@\���8���\����Fg��T6[ӛB��<"�Uq.J���/�U5��@�Y����߭Wz�V�����h�^��a�یYs�	FYCs��*��f�%rrO��G�ԫ��I�Gs'a��oq�CV#�D:�L�#3���2*@f[	�t=�r��o}�9��p����*��uf�1J�Ǝ��X��̈́eOE��T�.Dr\�1f nI��%�I�,##�M���Z���!�@�x�M�zS�����!���4E��U�r}12���Q~*�~F�VD���5,6������#���#�̕5��p2�p�^��'�ژh0i��nu�v����9Q����o:�~&63��?6����ܧw�d�q��5���'vT�j�<��Sxe�uҟ]f#���j����שr΁�y[���:1����Ǭ
��v����Q�9W*�5S4E�]��7s2
1̵��܁ ��
��X� >4�7KHu)�%��]�q�+'��#l�b�ׄ�����dMOd*��E%��.R_� �)����ZTV
8W���
��H��)�f�R_cJ��2s@�.Iʫ�-��66:ڲR��0@��Y�a���L}��Q�?G�D�/�| $=MB�H�N���7#���GA�٘o>d���֐N���Q]���#v�N���Q$����v���Xi+(�&��ѐ�Rfȭ�H�����W����{)�ȸ#"$���P���;��MxJ鷬�b�������c_��*�$%e9�MY�KO}��XI<��q���{V!4�
}����bN����P�e��d+0^�'B���5j�h�E��.�?p�!6&�ݕb�z.-K�S���(GYv��~i���u�{��)N$��0+� ��	l�a=q��-(�X���ќ���M�3'I�(p�Cn�t i;�N��2�
�����ȃ/w�O�ѿRo%-z�ş����9�p�8����t=��[��B8s(t�!ڰ���h��ި� �?0ߞ���'/GE(Ky�c9SIc���dj�i�����f�-�g���I^s�)�z<9�=��K�%��6Ѿ���5�,:]�U�U�x4�G�	Ά�e�l	r���S[SĳQw�4�~�����iEg0=�7�w���3��m��mwm�|�0�nK�� Wض��/�8l�N�y��u��3�P��Mp�н�� ���ˌ���m��t�F`ιxHʑ�7���yԾ^�.tgJ�R*RމD|/�s��A�A�)8T�t-�J�u�-�C(�7����jJ�S�1���f�[�pb#��}�s[���Q}H�MM�U:*��ߏ���$я8�Y8��U�Ζ�8?����e�i���ѽv�C|�A�R���B �4W&B�#� K}���E��-V|����J֑e�4aA�%�|�`M����R��(��S\��f��h��E�!%,�\��b�QdQH��$T������H
�ު�h,$M��Y,�m���3de|���6 ��d ( ]�pT�0_�tz/K|���fL��|��t�wl���_;U0u�a��o����%���$i�\f\�#��L,��|�_s�;Ρ�/�1.�ΜX��o�}���k��T��~��2��<&<��c��e3�����DJ?W�U����q���҂�!u
�Q�b��Ð�����A�lF_T�`�Tx��{o� �����F�'�Xl����K��ȎF�dk͋�W�
��	K��뚪q��C�������������G��_�"^�z�j�+���D�h�N��������>R�v�pBЩM_ k8�>g�hQ"�;n�	cfgz�o3��u�Sp�Z��\���%d@��2�9s����Ԫb�i�E_�Ҁ56��؟" ��`\-s��>}���5Ͻ��tU��������!��lC��-5��8����QZ.ĉ]��O��-�Hm[=��ss�������ggJ&*����I��U�X��e��H����Y�氍䃻E�:�d��لPC���3�(�of��x?72���{���ǒ�17 �>V�-0��)��.��SL���
��L�l@	�H���K�=U��`<���SC�_�e��-�6��c�/��Cw�g�g4��A�s���7ՠ���`Ȝ��!�2����h��Z��> �\p��gR���fd؁>�l5w��-`�~<d�$����<�˵�d�eVb���ℙH������aLQ4����c�hR��C��o��تƹ�:�g��i�#K2)�\<M�hvW�|�&u��;_W�a7A����Ǆ^�	�x��o��S7��-�|~���$�-h����E̽���)�ORH%�9͈g��G�=�h�g�M�:#%cx��&��,/h���ܓ��&c�N[7},k��a�o�EҴ���\����eقr�3م��2+�6��账����q��WD�h�>}-�B6�}�<@(��w.�o�o�