library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Color_LUT is
  port (count   : in unsigned(7 downto 0);
        switch  : in std_logic;
        VGA_RGB : out unsigned(29 downto 0));
end Color_LUT;

architecture imp of Color_LUT is
signal index	: unsigned(6 downto 0);

type rom_type is array (0 to 127) of unsigned (29 downto 0);
constant CLUT1 : rom_type :=
  (
"111111111100000000000000000000",
"111101111100000000000000000000", 
"111011111100000000000000000000",
"111001111100000000000000000000",
"110111111100000000000000000000",
"110101111100000000000000000000", 
"110011111100000000000000000000",
"110001111100000000000000000000",
"101111111100000000000000000000",
"101101111100000000000000000000", 
"101011111100000000000000000000",
"101001111100000000000000000000",
"100111111100000000000000000000",
"100101111100000000000000000000", 
"100011111100000000000000000000",
"100001111100000000000000000000",
"011111111100000000000000000000",
"011101111100000000000000000000", 
"011011111100000000000000000000",
"011001111100000000000000000000",
"010111111100000000000000000000",
"010101111100000000000000000000", 
"010011111100000000000000000000",
"010001111100000000000000000000",
"001111111100000000000000000000",
"001101111100000000000000000000", 
"001011111100000000000000000000",
"001001111100000000000000000000",
"000111111100000000000000000000",
"000101111100000000000000000000", 
"000011111100000000000000000000",
"000001111100000000000000000000",
"000000111100000000000000000000",
"000000011100000000000000000000", 
"000000001100000000000000000000", 
"000000000100000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"111111111100000000000000000000",
"111101111100000000000000000000", 
"111011111100000000000000000000",
"111001111100000000000000000000",
"110111111100000000000000000000",
"110101111100000000000000000000", 
"110011111100000000000000000000",
"110001111100000000000000000000",
"101111111100000000000000000000",
"101101111100000000000000000000", 
"101011111100000000000000000000",
"101001111100000000000000000000",
"100111111100000000000000000000",
"100101111100000000000000000000", 
"100011111100000000000000000000",
"100001111100000000000000000000",
"011111111100000000000000000000",
"011101111100000000000000000000", 
"011011111100000000000000000000",
"011001111100000000000000000000",
"010111111100000000000000000000",
"010101111100000000000000000000", 
"010011111100000000000000000000",
"010001111100000000000000000000",
"001111111100000000000000000000",
"001101111100000000000000000000", 
"001011111100000000000000000000",
"001001111100000000000000000000",
"000111111100000000000000000000",
"000101111100000000000000000000", 
"000011111100000000000000000000",
"000001111100000000000000000000",
"000000111100000000000000000000",
"000000011100000000000000000000", 
"000000001100000000000000000000", 
"000000000100000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000"
);

constant CLUT2 : rom_type :=
(
"111111111100000000000000000000",
"101111111100000000000000000000",
"101011111100000000000000000000",
"101010111100000000000000000000",
"101010101100000000000000000000",
"101010101000000000000000000000",
"101010100000000000000000000000",
"101010000000000000000000000000",
"101000000000000000000000000000",
"100000000000000000000000000000",
"011111111100000000000000000000",
"010111111100000000000000000000",
"010101111100000000000000000000",
"010101011100000000000000000000",
"010101010100000000000000000000",
"010101010000000000000000000000",
"010101000000000000000000000000",
"010100000000000000000000000000",
"010000000000000000000000000000",
"001111111100000000000000000000",
"001011111100000000000000000000",
"000000000011111111110000000000",
"000000000010111111110000000000",
"000000000010101111110000000000",
"000000000010101011110000000000",
"000000000010101010110000000000",
"000000000010101010100000000000",
"000000000010101010000000000000",
"000000000010101000000000000000",
"000000000010100000000000000000",
"000000000010000000000000000000",
"000000000001111111110000000000",
"000000000001011111110000000000",
"000000000001010111110000000000",
"000000000001010101110000000000",
"000000000001010101010000000000",
"000000000001010101000000000000",
"000000000001010100000000000000",
"000000000001010000000000000000",
"000000000001000000000000000000",
"000000000000111111110000000000",
"000000000000101111110000000000",
"000000000000000000001111111111",
"000000000000000000001011111111",
"000000000000000000001010111111",
"000000000000000000001010101111",
"000000000000000000001010101011",
"000000000000000000001010101010",
"000000000000000000001010101000",
"000000000000000000001010100000",
"000000000000000000001010000000",
"000000000000000000001000000000",
"000000000000000000000111111111",
"000000000000000000000101111111",
"000000000000000000000101011111",
"000000000000000000000101010111",
"000000000000000000000101010101",
"000000000000000000000101010100",
"000000000000000000000101010000",
"000000000000000000000101000000",
"000000000000000000000100000000",
"000000000000000000000011111111",
"000000000000000000000010111111",
"000000000000000000000000000000",
"111111111100000000000000000000",
"101111111100000000000000000000",
"101011111100000000000000000000",
"101010111100000000000000000000",
"101010101100000000000000000000",
"101010101000000000000000000000",
"101010100000000000000000000000",
"101010000000000000000000000000",
"101000000000000000000000000000",
"100000000000000000000000000000",
"011111111100000000000000000000",
"010111111100000000000000000000",
"010101111100000000000000000000",
"010101011100000000000000000000",
"010101010100000000000000000000",
"010101010000000000000000000000",
"010101000000000000000000000000",
"010100000000000000000000000000",
"010000000000000000000000000000",
"001111111100000000000000000000",
"001011111100000000000000000000",
"000000000011111111110000000000",
"000000000010111111110000000000",
"000000000010101111110000000000",
"000000000010101011110000000000",
"000000000010101010110000000000",
"000000000010101010100000000000",
"000000000010101010000000000000",
"000000000010101000000000000000",
"000000000010100000000000000000",
"000000000010000000000000000000",
"000000000001111111110000000000",
"000000000001011111110000000000",
"000000000001010111110000000000",
"000000000001010101110000000000",
"000000000001010101010000000000",
"000000000001010101000000000000",
"000000000001010100000000000000",
"000000000001010000000000000000",
"000000000001000000000000000000",
"000000000000111111110000000000",
"000000000000101111110000000000",
"000000000000000000001111111111",
"000000000000000000001011111111",
"000000000000000000001010111111",
"000000000000000000001010101111",
"000000000000000000001010101011",
"000000000000000000001010101010",
"000000000000000000001010101000",
"000000000000000000001010100000",
"000000000000000000001010000000",
"000000000000000000001000000000",
"000000000000000000000111111111",
"000000000000000000000101111111",
"000000000000000000000101011111",
"000000000000000000000101010111",
"000000000000000000000101010101",
"000000000000000000000101010100",
"000000000000000000000101010000",
"000000000000000000000101000000",
"000000000000000000000100000000",
"000000000000000000000011111111",
"000000000000000000000010111111",
"000000000000000000000000000000"
);

begin
	index	<= count(6 downto 0);
	with switch select VGA_RGB <=
	CLUT1(to_integer(index)) when '0',
	CLUT2(to_integer(index)) when '1';
	--VGA_RGB <= CLUT(to_integer(index));
end imp;