library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Color_LUT is
  port (count   : in unsigned(7 downto 0);
        VGA_RGB : out unsigned(29 downto 0));
  end Color_LUT;

architecture imp of Color_LUT is
signal index	: unsigned(5 downto 0);

type rom_type is array (0 to 63) of unsigned (29 downto 0);
constant CLUT : rom_type :=
  (
"111111111100000000000000000000",
"111101111100000000000000000000", 
"111011111100000000000000000000",
"111001111100000000000000000000",
"110111111100000000000000000000",
"110101111100000000000000000000", 
"110011111100000000000000000000",
"110001111100000000000000000000",
"101111111100000000000000000000",
"101101111100000000000000000000", 
"101011111100000000000000000000",
"101001111100000000000000000000",
"100111111100000000000000000000",
"100101111100000000000000000000", 
"100011111100000000000000000000",
"100001111100000000000000000000",
"011111111100000000000000000000",
"011101111100000000000000000000", 
"011011111100000000000000000000",
"011001111100000000000000000000",
"010111111100000000000000000000",
"010101111100000000000000000000", 
"010011111100000000000000000000",
"010001111100000000000000000000",
"001111111100000000000000000000",
"001101111100000000000000000000", 
"001011111100000000000000000000",
"001001111100000000000000000000",
"000111111100000000000000000000",
"000101111100000000000000000000", 
"000011111100000000000000000000",
"000001111100000000000000000000",
"000000111100000000000000000000",
"000000011100000000000000000000", 
"000000001100000000000000000000", 
"000000000100000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000",
"000000000000000000000000000000",
"000000000000000000000000000000", 
"000000000000000000000000000000", 
"000000000000000000000000000000"

);

begin
index	<= count(6) & count(4 downto 0);
VGA_RGB <= CLUT(to_integer(index));
end imp;