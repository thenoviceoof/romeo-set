��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�ϗ7�#���H�����u�g[iˬ���t|�3���ҥ�ys�B�@Yq�"F}�\"QY����#�ڇ7�\ӷ��繟��1W�k���q�u ���{�m)RM�S|@�����ͣz��yʿG��O�Yg>�s$h_!��-~���=wx�=�M�����/�mb�K#�� ��1��W�i�{,?�EM�N�0�K
䧣�:39ok^�(��-���V�f���Sk�	����}ؖŸ�*����~������6l@ޱ����t����_.��±7�Eۨ[�ܐb\T�8�����"��!'���^C�he�K�Zw��J�;��E���a�BnB��lje8�i�U��^w�K�@ܚ��^<'�������������a}��a��W��S��!�P�:�ޓ��|=ǎO�k�σf&�_ K(yǦ�+F{v5�X�x!}e�y�D��"љn3]��6:�Ѳ=&:_��h�,�klf�es�4�=|��-�#3��r�E8m>�e7�{�~w���O3��{	 X�n���7��[��{d�mҫFG�6�ݝZ���4́���GF��yw�D��Օ��挹O����[�K6���L���ڹ�\Z'�
���lS}d}��w7�� ^$�j_��묡X<P�`��&X���xRq�y��G���R��B�}[�b50t��j�k\��Ju�a�V�ؒ���w�\%RF�Z�購�:*EO�GT+���,��B�/�9K�5J���t	���y"q��yǕR�<�]���>{�t�f�'z�(*��l�����'J|N�]�F����Yz�ȅy��/��)�B��
�vu`o9M5|�Z�e������gM"���C�W��f,�o�`��<��Xk�:�s#�T��/q�PC���k�!}5������j��b%׊a1-�b��\%猢��S������Ew�Z���UYwds�i��;�IT'q��z9}j��!/m�n��4�Z������ء�\��0d��>�fZ{�>�Q���}o�x�/=̪Y�I�s<T�y-���G���_�җ���2���5�g�$K�+�'y��wj�%��� ����s�ٸe�p{��V�$C����FQTX5��)w�"��c��Lg+Z�fvV@4�ZP�>l���
�U��������tAĪj�k��V����>lv�C�/8��M�jR0�:q����Tԅg%�L�:�����t}W�/vF�XȰu���*_=�Ҧ�/W �W�J��k2|�v����Q�o�2�l� �@��n�S&E����q;�Ǹ�(�b�?��&�pAM�� k;Eb���7��U�U�k�и}8�+9$��'����ݧa#{�~P�C@�u`�#����]�S�N{"C=l
�i��+*<�L�n�k��STA��s�%�X;�y��@����L����n��e���-�4���=���t�X�	���B�`�K�C���Ɍb��8!5te���i� �������9�E�y�w��ܺZz�
�5�_�w�.W%x���|�	
�Z�� /��x���f�-H>��|�)O�(�x��:E��&��Ͳ�Q����<>�E������B����
\�t΍��9��Ȟ��\���$�z`�� �1n@4/��e�P��$���u-��?�J�$?���Q�Mʕ��[��y��ن@0ha,��t�H���OD0�p�{O��M=f~-�G����(*��!m�Es'�#�A~�G���yk"�ї�����!A.���Qձ�&Yeis?ޖ`r4��9��7H�͚J9i�Ň�yʣ]��,�y��)�Wz1����?����Wt����� ���� �mT��"�\<��o�����D���^ϝe�x鞾�F̂���ˁ��ͪ΢:yz���Jc
��CN�!=�,�]$a�����Ù���2���rTc���Z�=HZ�$�Z��^T�{)�ȧ���_ׇ߹k ݧ �dظ�z����*����D��٥=ɬWb�	օ�����^���Ar�pLPH�7��G(�.O�]\��Snf�ǯy��(za:e�^������.�Ƭ�r}�GMP�s �Ǭ�����O�x����Y�T��3��`��3h�s:����\2�d�;n-�q8���FW��>3�|o�
|�ÿ��F4I����[Lb�8��9'�Yj�l���[T��i�V��p���eƤ��h�9���`=����[Pf��c���#����4�7����Y.@�ݧ��{��Q�MDm��D������C��2��]�4���vK��B����s�6'.s;�Z�U�e9J�:9�7��@T�_��ꐜ�M�x��>�`�� ���"�k�(V�я�����5��GS����ׂk�M���I	ǳS��Q�N��P�ĜF�GA���Wy�j-���D�k�*��M����ՒJ	�q���Y۩>q�S���R�(Em�F��\���-�h���Pj	M4oı����DN�����(,�,�|��SO!A�5��.��2�ɉz�	�K���q�'�=[ʭ|LX��Q�h;vn�S;̝�Є�%/o�f?*���[�B*�z��K4��)�D�gz��+.ݕ��c��%�V{X,,7+M�0cc��;L�W���zo��ϖQ���"�L7�k��1�鲾ě@�uo#]��` �00�v�3)��e�o�g9Д�(�e�$��5�z�m�7*'��
�.�J��ly�L:,ۨWu0B٤����?��RĘB+%yY�|�Q@������¯C>�<卓���<X�dI���I:�!�r�4+#(lpؒ&1���эb_�+V"������a!!�h4�B��PS@ {4�i.����eG�\�w9v��<��pp풥�OYY�0������Co�gFFp�[�|o�s��u��-W/�Hx�o3p�+F�;Lг6]6b��$�^W(�,ބ$���(�?�g&kyt_�e���s5���VE����{l8ݎ��Z�x�'8�^+��Wl8˧N�]v�Xѡ�t �m\K ���a����)\�$J{�[�=�4��h�}�iy2Z��TDy2@��k�N0��~���qt�x)�{��N<��LW`��uT�*���(�;�)��)���@N{��'zoT)G� B|e�eH\�(8���@�,�V�6����r��_8K�E:��&w �aeC�&f.f\*������2�e��C����<���
0�?��u\kYA^M��*��i^�X	��0]Zs��))�z	��l��8k�aNe2��i��3V5��]��zv��� f�\��$��Oƺ����Ni.�q-�Ӭ#��X�	O6�<�)��c�Xͱ�3��X�Qw���8RJ�x�(��xsC�-�
;Տ����px��'lHR
��Z��{|�{�1,
 �e7ų��	f��������~�GPV�S5U��0���(�ẗx4��������W��H;�*����j�;��������f�������D�Q�H�Nڡ��gT�Aw75��7�:�C�X��4�>�<%�i�Z;n5�VJU}!�0��zu3���ky��`0��M��
��j����eqw��T�xvB�c�1EzhMP]0X�X
"4p@HHW$�ik\9��D�{����i��Ԉ<�2M�v���,�@-q�%v2���,�=��埱�lѕ#��
%Z˓u��O�
�q�:0m����K�Pu�!0�;���j�\�Kyv�k[�0z�GN����ժ��R�Y8-&����i�]d���� ǹҷ��c�&�qO�&o.F�Eg�=A#%0`�Jn��U5�I!�d�l�J�J���V2Ylie�K��:_BĘ���;�����.B�|d��`�g�- {�y�Jl��L��&r�6 x�M"�p{�[�{Wc�=�!�ٓ.ۓۋ_��I[n^�� L^�
��2���I�R@쒬���H�n}��ఉ�y�fÅ	���>�,r�-�-^�<1�L��$��h˰���L��X�ibI/�K�J��jXc�n��w<�A�J��ȅ?����N�ݤ�z��5H���ߺ�=x��S�ˉVH�x���Ր����p��O(#	�ӽݸ�� '���⩊<0�v�o����V*��Kr-�I
�w		Ŗ��i��|����9|��N�3�
(=��0Sh�@˔��f��Un�6�V5Վx����o��B<�99?P.��/ H����gY#0�<	��� ��+PZ�E�V��)�J
��s���.�N�ΙyŽV���_I��O,��`�'��<|��YЗ�[�QҨZe�T��B�0\�R�:�&�>�B�Nݠ�,ʝ����/��� u�=A����#��d�
z�U�x�5����T��4�sK���m��E5�rfcg9bx���ʶN��V!�Y������)#-D�+)��9D�$���+iV�9�SaP�	�p�~>r�o���n17�7RRZA77e�)*D���˄ߣ�d�f��������)�%��< J�v��)4nO�D�Q�)�wDX5�@a��=�;�7��a_w�OR�zw�r睟�;1�?���17�0F4OaQ���܎��Fk��bp�k��o{��u�������?z��dl�+�H[m��5��xg�#3&4}����J4�
(U��Q�-���3x�T&4H��(����|"��Z.��
���hN���Llk~n�q�A��1��x��Gޓ����bt$���pԸ�P��K4Ķp����w�Kf,8{k�dA�i�p7��֩�i�~}�G�d�Jn/��1?>�n,�i~�n�sh��D���g)O5X��u$+�f���V�z���\(xL՝\�GaIrE/`;�&���m.�7
�\��y4�Ie^S��/u���V1���?���B�e[ '��{��SB� *6���k��� KR����z�����h��g�x�ǭ�ʧ�Č����J;)s'W=w���z�9Ich)=�_�#8�{���\����=�/�`/����ԂapQ�����X�+�^j���`0H�t^͋�Z���u�R�Nl)$�^�w�*<�xG����.����Y���Qp�wu�y`����R�Zj��@�ery���y��	ܠ���w���$�]u`1�f���pd]ӏj��u��&�fU��¤��7��K�>^FA@gp�
��J��N�l��[P��k�Q�����Fy���Un#g	��g��'�mO*��P���N���1�>W��c��l����Nֈ�=��k���6�fsm;�\o��m$hjAW~$��a��o��`�@�c�=7»9u�{^��%�ؤv�F|{c�;ǉ+ac B�f�R�3�g�S��J�Z8�)р���F�OA'y�[��⫖%
�L �0�}żА�f���,^���kи�>l���Hf����j��G%�=�ܣr����dYD}q �y��Hf�
x����F���8#�B�R����s�[�m�Ow�C��"���F)�ޜ6iP��k��ӹ�z����T�;�o�Q���×HE���n� ���z�f��?:N�s��(�j��W*s��u�f8}�U�K5�#a�5+��V�bKI�R�K�rQ�a|�U]��xq�����n���]&%�\�/�a^�:�3Jkc�'l�n��ǎ�5(0Hש-�u��J�z{���@�1Wӆ�̀��������VCQ	K%kl�b.�<�Sx����c�Ü�B�w�1ڙb;u��Ʊ�������50X�hr2�G:�����JI�'�IO�V;Q)+�V���.��wh��.4*�gH:	�(7-��[X�DT�L���j,ӏ[���e8�'xd�O���*���Yrnx(������x&,K�<���d�SU�ߗ��J	�7��J?H�ڒ�@�f�p�"ћT�#%�E/}�K����>:E�����k�R.��Q/��7���%�ʪ�b��|�/1�b���谕�TS���~���*�5GKf�/qk����F��TkF'��ReY�KmVv/����-B2 �`��j$����M�FGC�`Y����EB�I�e����P]N/:��9�_�����N.��s��s���4]�aI�5�
�l��N�M��5����W�!�]f[���h1Ħ	��Ń�_ZX�l�է賁�U^Y�E2|��lƉ��^[)�G�����8�%2�0X�D�t��¿?B�O�7���ū̠�8�N�"8�;-�j!����Wk�}/����ȳr�6�(�e�}T��2�U�P+@ސ�ӆ���AϮ�R7D�D�/+��oC�1�U�#�i��_p�4�3��G%�]#��NwN�zY��Vۧth���������TL�`�3g�;�e�a�@L?���t�mOWX�p�s:�V����a�����C�!_�I�w�)���a�������xُ�+����R ��(T�ierUc�4���t+!��cO0=n��+�CDp�!}g0��I���jH �A;:.4bYv��#�w�O���c9�@	�K�5���Z��
�$.��c�+���cr�3d��$Ч��ˬ$�G�-��n�%L������Fdi2������t�H�y�,���v �$�=Ͻ���9��[��r��5��9�J>��T,��X����ʟ��EQ��)|,��C�]8�����y|dާ*��D~����#Un+~.�$�x#b��v4����v�=�Ohيr_���1敾W�	������p��1�t�.4æ�e4~��"8/V������|*������贼�((@��]{Z��H�� ���\�s�w�G���q't����[!`t,wNV�8㾽�-_q3��hD�6H���%fv-��4���a8��5�N:�)�[���_l��F�yXX�������+��x&`,��Z�`��7?g�/b�ɀ �9����/���o.1Ʒv4k=��z����Xn���0�Y�4!���A�!���mK�{��FE��Ww8��qeVd(�%J¹���0��ܹ��;L#0ݱ=���]P�j��"]��i�CC�&�GZ�VY�+#C�a�@E@���2�� -"'�xf��s��6�mY2.	��P/�G��$s|��AU.�M=��+p«3TF�Y�@t,�Qb
��5�Xj|�*8��n4�]��ii�l��Y6,c��1\���&�����k���e1�m�<������T�=:�#��Uy:2�� a�C6�0�gܛ�q,Ix����Z����-�e�JB� jnJ`��~�1�q��ڀ���2�j�Q:�@?b��1��;��,x&b '�8?�`S#��B����&��iB�]@�L�#�/o[�oI�
�:�4��o�ͬ)�K���@��
Nf<$���m/!�"�׏��3� �����T��Ƒ��=��y�-�r�1! ��1ix_����v�3BR7���I�]��)PS�ҧ��f_kA����Q?m�������hc���P�z%��,~k���w�Ͷ��Ξa�Q��ܪr/�t�EuP���6�f�������a�����W_�J@KL�9�`�#��-疩/bl�FW!1�����*�����wZ�)��f���ԃ��J�A�.�h�@C'�����*�T�~��"=��rL' �vC���I�{�- ���&!K(�.�s�����P-��4�Fo���E��w�s� ⢽]���-\O'�߹d�U�	�jH��ԝf4�;rG*D�_6������~P!Z?�;wА�T�T8]�_�>�)M�����tXz=�{���4��rץ(i]�v��Lhϟ�fś!Y�K��m#�/���~�J�	����*�o#\�H�!>3}-����Nl��M�m�__o�`���R�5���R�e���'5Q�Yo����Ø��ԡH��U��t2�o�	�		�*��c�lxe �WEmK��z2��347Ԛi���䩰��bl�Y~��f��Wؾs�ڝ�&Ϳ�	���~'k�gC'���&7K� ���œ9!�;�Ш�"�9����SrEƷ�������Wo0�f%l"�A�M������Nx�9�~#�-Oy�e������Yʛ�=P�[\�o���)ga.�� C��߶gk	w\���w9~l��z5Y�ڻ(�`��,�U����<����kd<"�Fk����i 2�*߻�����m�i����*`��Zɕ��:+�5R/�,M�lb�O��.�� �s��ۓ�e���sY�j�w�P�ku�bm�D|�G'���I�;{���n��&�&��{��4fk+�[���0#��u��%�YǷ���D���ޜꤲ\yjK��~Ɯ��1l���
������i49��\odf��'����$�ۤH;�R���}	]G���T��uZZ�{@ߒOzQ�TY����!�z����ī�jL�n��m����4�sEu�Q�-�	�,5ёZ��C�*uɇ��?'�G�;Ek���ʣ�[��f�;l*�д�#�斡�{��߂��=���"�z��KR��r8]��D7X(�ﴥ��"K��$��|Ao&��v�����75jV,Nh\dΞ�� �I�%h-��C���Yy�1q*j���qN��~������]gG�L�m"k>�����:\���٦' �O\����E���׊���;��;^&ժ�k�P@�·3�z�eȲ-�N \�|�}"�h�e0�����'M�`�x�R�U�"��6�ܳ��ou�ȋ%C��������I�<R��������N�@��J�ٶ�٬�u>;����x��ýCۦ�25�N�S6� �dS�b�y������c���U>Y[|����W�D�;c)f���YY��ELtN]�wg]���.T�c }�f��$tեn�����Y?W�NO��8�w+~]_�*���2�x�e�bq���F��	��bp�$��=5-譖I-3��Bj�?"!�v���A�Q��	��%��c{>o��!�Vޤ����j����b`�P�w}� �dJs)׍Ci�Ej��$��wk���\�
����.8ɲTݑ�^�h��L��?�F��a.dZZ�d�f'gF�7d^ h�ۈ0�I�汓�=�|��^kla+�O���N
�+�S�>zxM��d��U�P��{C�L�Bv�v4̿����q���\��k�G\)/ Q砷D�ǌ}��I���1�&�����ZtN�*�H>d	�3l�V�@��`]����Q��YU��1�#K��?N&�=5��|��ž�%1&���u�)�T�ڞ��p}8��o�����y#�)�����5�5:�'�ũQי&�'��5h��{ֈ��|Q��8
�i �'Om��CK�w��=Vlos�n���a4H&+ؕ�n�{g�|VW�W���LÌ\�Ne%΄�X��h/b-�k	�joz�.�Sn�k��!Ƭ��6���Z����5�;��x@�~Q�˙�ɿ%��='�3�{#���{jᚱ���r�f`��_��+5�&Q����� +M�/���g�@�񡰧�Q�̽U��ꜿC���;��T]�a%S����y�e�e����5:	����b�m�.��Z�5�;;�a��EZE�o�N� iީt�������V^7d�pr���Rʉ5�R����W�5C	�R�y�y<(�wH�o?����.�Qp�DK�}&HG��38\h��/o�\��w<h���Dd;_�cїlX��D�^$/�ۭ̐ߠ��E��?��j�Yz��OE¡՟!U��@S}�G4zj�m=tr��0����ۼ H
�hՄ�OZM��B+���S�(��<��E��>�J�5D�k�0otN�T��Q��Gh�6���^ѷ����3��p#j/�O���� 7���n؈QXܢ���w�u��c�AX�^O~��'^�I3h]�����4sώL!Vr�7��	�g<8a���$i;�
�{0�p*�}�vv��#q�9y}֎6b���l'�Ә�D�Y�EfX�@������5p�����s~�������c�?�4��Y����?��*�s�PK2 �x���x���w��)���X��\��f��K��""�Cx���y�$~�BRvݧY������*�xUhnrY*��Z�U!�%X{�
��T�F�H^툉��s�
ncX�춼�7��\��w�v��$�T�)��w����yp����ICXuu��H�f�:�ִ���<�*Ӭ����9���
���B�ž _�ݥ����HH(C^�#-;��KZ�%�ǐ�D>���?���-9�9<Ԥ��u����_��E�[ꇘa5/Ia�f ����"z^��}H�`첒-�k�)�u:٬9�8U�6�ݎ�~A�E���D��z�h���S��b�W���A��n����*A�%�sf^ �2+�{�by��uַ�#xt�~���*� eT����N�d�����ms��+c���
[�*q�s�*��d,�b�M����͕��7�h���e���{=#�����]��0�I�q8n��h<�P����Q�O���,@4/lS�PZ�ar�&����ƕ�X�=��-P<����&�c^��d��;�`��Ve�^�5����'"'؅�X)(S&�z���J��<�vT��`�'�q�Q�a��%��6Ϳx0��hȡ�pO *u�-��Q��	?C����u����E�C���O{R>�;�Vo��]�J�~��5�:f~. ��r��ͥ|s��9T#A�g����.�����~r������96�7SROT��R��g ��KԞw���G7ߣ�6�u�tn:&��6��|l����K"�(�&�|� K�'���{|f���-ؚWy!��8��?۹�K�\�U���b	��v
�l�������WWh���x�H�����es��b���#!{%����*�-}�{NwK��RۿiX/�Z͜p1�o��nma��-0���;+��t�a�j��4Մ��i4�i��X�rp"���W����S��d椗���%�?�g/�9�c�p��x�4�w
�7@Gpr�P������o��epvRK���J��Ҥ?r����''x+s	|m��;�v���> ���IYH겆���6k���L�O���3 �^a�%y��P��+;��u��yg�`��+k\�������p�=*y�j��r�
��C#�<�^r����V�dv�r��X����!����сj-�[���.�./��T���;^����/A���0�r����3����q#��e+��V��E�L��~� ��h���}��H�]{&k>*��l0�Ne#�b�)�ҕ�8	A]�{썌��*�ʠ<�.K�fVe�fS��*63�5Ӟy�4��?�R�9ǟj�1��_���Cb ���PF4��@T8�e�����1߲H��W��gY{���)�����і+ח�lgk2�������6wq���)��v.����Y��Q� �>	�&q�`�����S������g�e��&����&6^ོ���ir�.(����r6uJbF��\oGo�
�bE1P��/�;M��6-a|�A��T�('Q!
�T�v-�S!�̈́_�9��b9->oM|c"�Y\Tn����df��+�*����-�:ni��jM�7座_��B�^�u"ͩ ��%4�s�I�s�z������z��c[�4��˦��7����+�`���S���#g�~�`�@:�s1�g2�p���[���k�$�V�ɲ+x<h&�#��fp2�A�A�7]����Y�W/%G�I�1W
��\�s.�Tu�t~kdW��~�-����Mh����=ܟl��QV�51�SX�,�]�fHWU9�h���oa�՚ ���
J��t�!�;H��~}i7�<�t�0c%D�>��q&;x�F�d�f�n�
�w�Iȯ��i7D�R� 3�p&�%��F�m>�E+n��FI�eϒ��GT�8F]?�e���rV�"�6I�W'ĉ�&dMP�B�5���5��:~��A�=j�2F�(Ø-�կ�?�|e�#2��W�nE���I���C���Q,�oe�շ�)b�!B^�h�km���L���(>���Nk��ۉ�b�Z�/e�TE2�Ͳe��6`dv8��k�����Q��j��Ks�E��q�W�Uc�"�XYz�w%%#쬏6Tx�����
���L�� $��>�;�ѻ�������ϧoe*���S�"�ǩ�E��y�8$
P7!,�E�����
�!+�Q9�c�*�@o�D�L�߫Q�Es�M���<�n��7�F�t��A0kI�Pg5����0!ͦp~i1�lՉ��C� !w< �� �}�����o���v�ҏC(;������`4wϪ^��An��m0�� �=?:1���e�-�9�mՄ�CL��g�e9�>Bv/82,�xgS	���@ ��Ly�,�����;�L'bzϦn!�g�wG^�f,c�N�/��	��N<@�k�.s�\���B�~�7�)c�GM6J�qW�]j޽�Y��Vn�ږη=yL����o�]�S6ĺX��c/a���(��.�t]т�_P�G�<c]��/�L� ?�����"���N�upwMٔ+	��fD��N��e�L˥m.��`�9Z�۰C42�_
J��B/��v�XU��L����^r�uv�r֪�-Z��v4����)r�ۣ�:4�����?\��eD�6"�4�̠-�����!V�Ug��y�9r�ujpXϽ��a�sP.h�JS��T�]��B��v�r�.ѕ?��m�'O��j�S9̌v���4������6�X�8׌��H�"p6yYF�q<�����Oׄ+��nZo��h�!�[.��b�E����`E��K6��n(N�n튱���2�P���c�'��������V n�
�]>�e��˓����O���fP�nN�Vgc���w���h�QBm�W�N��T�Z�wCX�����W�#I��W�Z�i���^�,.W��(A�C�*A�,#�>aϵa!�L>ۅG;f�=+*(����]����ϫRV�Ƭ�Ǟq{�gY�������<! d���+3�>��[�)m?��N��z�QLZ[[(M��w�ʱ�\�6�b"�޹|1Ȼ���FV���T�DID�p$+aoc�P:�t͉n�����a� 2�G�ż�����O9�=��I���T�1�S�Žp���rZ�0Q��NK7�2���N��vD�ێ�z��$2z�T�F�b��@�@o�;�I]��y���=�3�_������yd~;"�<����Y��P z�b��8Y��l7>���ϧ{�(+�q�Y/~Xt����$�.��{Ǌ۲F��m�4%Ѯ�����*	@U�"���?j֞Y�+V;|��VH���T���d*���S~k����_>��������#e�	wC_1�&�ў�!���~͹���[�k��2h��{h�UwW�>|:0�nȈ�FGe͒�%��'�����e|����b�]F7�Np,r����5Fd�!2|?�����`�i>VMT��X1)E�������p�c��*��\rfݽ�c�QsmY��J6	�q�׋V�fK%r���h��ћ���ޣI;�b@A�S+�Rqb����o_"C�������W�J�/����59t��Gd������b�<&�9�ߤ�$�N��5Z}�����U���W1�ӽ.~�3
?t"���H����T�s|��Y6�d�����N�q���bN����D��ŖL%��b���>�T�ٽ�4%<C�>W��f��`s#^���@I��dl-|�׼��0��&��K=*�G�C�kX��T2�k�RMI��Z|�����ݍ�j����6T3�����^f�p� ����~�U���:7;�f�S'ep��^�N�D�Bs�����k��%d�laB��O���*�����x㚶�wbj~�G7a���� ��)I�?,?3р�%U(M���%��6��!$e�"�:sUX;^2=�x�h��frș�����>	e�~]�U�1���\�:�2R���A;]�%�*o��:���N��Zy�T�����`�=?���Sq��JW�O		{�- w/#�S�H�P��/C����?R3|���й�zmO[똿dkfS�!�޳<g�V�a����t�N�V-� �eȪX%b�(�)#DoN}T�xNW��52Ӭ�܉�J�-���3��'���r]�DyGC&�����n��Hk�9O�[��#�����̣�%�w�C�+x�pi>S�ȑ����������~�'��+��Cv�m��IX�)n��R�"����Ƶ�S���)]G����[����IF��Ѿ
L̺�Ke�J��,�i�APV������K����a����D}h����S0EAKTCK�]��j��?�sd��A<C	åCW���NE��6	aΛ���./>��k񊯚p���&�?G�sO!,>W{��v��w=��ZJSz!*3��1*��Q���҃�0�ڐQ��m�Hΐ�3-�Mx��\�G�eQy~��#X�4ϟV��%YH�7a�0�7P�\`Q?��5V<E�*�xН��r�Z��[9nv��Z�Fb���e��8�hd�����+;:P��	�'�O����J/�e����ޮP��w�t>��k��	�����=��ɞ�*��H;`��Ǹ�*J���b�*0ko�7�W0^քىSKVzה+n�����F��tk�wh�e)Δ�m��ʝ
�Vv�k	�����
R�*3\<jm�P �pX�l��m�bڪ��J��^��������6wq��:"�TQ��(k��A�m�VlD�o�7g9�Ri.kD�����Q HdP�/p�Gw�PXTEB�&��/�dGCn�������u
�63��T��� �����{�f !;t���g������R�8�6�a��k����]��ܭѴN2�gt�6A?��YK-�$���@^}<��m9(��#�����cy!$o5:DC�ev�B����F0�'�s�1HG�	1o���Г�X����r��>��.�IPY���5�� ΃�8�\�A
��0:������_mbE�nM?C�J
����Dm��e7sAs��s�sfR]�!���F/�C�8�ܻ��)ҝ�?�s[C��x��TvBN�+.�J�ǋ��n��nkK;L,,�{L�i�i\}pB�T�B�S�}���-�M�*����0��#:�j˕! @��Me@�	9w3��`�a��ޯ���B#ߴoҵ�b~������Z� F,�ŅҾ��Ē����q��kJ���_�)��Vv�ת?
_t=�2t�1OoH��'(+l��^��`+��7��RΈ�0��7&U�o_?��'?�v�0���\O�!�<raa����n��"�_8�c�Ժ�u%~;��Q���kD��K�%V��E��^��_�W-��:lUđ���3,T{�V�Ou^/YK�x�gD��d��"3�HMkX�?�|��äje�=��;9��;��h#�f4���k�u(e���h����g�ȍ~�����e����᳸�hS�0�L�Ӵ
�R_��PE�b4�C{�99�ky*ɮ3��*���±�K���7�G�dv6��>��ہ�l�'�_cҌ�� 60��ZR�@n�j�m���꼙9+�5�*��E�h�'.�CC�6��f�|1�Ǒسp�oȬOL�N����.%�Fn�j�=cs����[���S܇��S��
��v����|��o:4i�
�X�<g],�{)�G�!��g�uV�3�ѩk���ٍ���D��]j���ғ
xL��;#�i}NxR߳��*5:I�Ȫ���� n1��gy�7��FW�tԩ�AՁ�wh�ěҬ� �"\k��#o��]���"��UP�3a]�,�ү�}@�I��RJ<�#�1����� ����դ�@o1#߻����ܠ�h}�o���3>�r�ks<�G�r��<�@�	#���
�����D�J�򘩴h�6��'��ȏ�sе��_Ri��%c�(��K�O"*AR3ϕ���)1�L z��l��~�Fu?���@Y I��<ʄ�a�'�͐����1@�|;���gw}�����X�7��)��1�9|�u\���-�4�^���	�A��]��m���l\�Nc�A�Ãg���uk��8⿈=��>�� �ܟ!EM���j����K�,��ߕ��"�,4��3�o, 3k���b諽sN�E~$6���>�b{��lɞ�����`��Z,���gB%�&lX���� ���E.��覸�ߘ_�e?&�]�� E�pS�˿Q#䔬���WUX!]�v���LIw&�,�7�u����ͯzU��6��Ȓ�[�'REd�\5Д�dϨH�H��, d7Rf�>�c�7�<o�\$<0ܪ���_9�h�q�IA�Y��*��o�l��eB�M�?̅���c4�D��PE��x�tDA����W��H�[D�ޥ���Q�>����\n8�z�!}���@�#n(�N�N�������\�ך���<���%���3��?m]�QM1bW�����d���xL��vnYs���;�n�:����,�P��TZ�e!��#�;t
��꤭��vf;� �=e+�&N��ߺ��QY�D:��-�p8v|I��N��˭�7i^ݱ>Vf���j���,�E�u��� {�N���pOVb:�2���czhl|��YpE��+�DG�����3��[#����*5�f�'�fl�d��YZ<ȧ�z�͸��q�3k���mg��!��!NC��/��9�����F�>w��Yғ9�={�l��,���Q��Ϛ���wޓҭgDP�����1�����V�1M-0��^�e��/�:�HZ��beQ#�(���ǧ�Π�i���f��垣��	�P{�B���9�('�"O@9qX��7�� �W�,�M� ����g5�I��r��Y������٤x�P�[��
&�h���ә�bU���;���HoHg�į(�W�c�#����`1�{�� �r�̺D#9{��<������"����Z&���r�>	����M<a��}}7xh.C����b[;k���3釮�mԓ��aL҅����ԯ%\������n�9v�F$9�56�n�dY�sq_SCOw�UY��?� ��T>��\����F�����tE�|������a��N}�}i��&3�Oz��AY7A�Ӕ�/���f~�&����2��N-�H;�(��IÙ�!t��Uؓ�{M���hM����e����ʙJ<�m����3;�H��
R�+̇
��??�̵?�ߒ�/��n�:]�9��h�� �O�p�l�V���E��^�]�mʨc#��+1j6p���S�"|G8#jf#�ԄD�R�F��x��d�;�ɭ����v5+�z����Nk���fZ-۶��H�6�O�J����V��[Ja�q��3��e��_�����"� �[�:��|��?D�D�[���=��|��:�0G],�B�t���n��M��v~̮��G`WnHY�i��О'\g?�! )ίR�k |㑶ё�9��<E����?��Or� 0�T~y ���i�Y�R/dy<Z����j�{U`(�W)ǴGv�RW~�ǅ"�Ѣ�*����R�e��n���M���^�Fo\7X����y���KN��Д�Z�
L.�7�a���ڟ4 O��G\
��{��7,�u��	z^S���O��I/�w)[���5�sZR���c�̚�C9ק�ք���ҡI4!��!��D��7�Ɂ����-�2�]䶙��Ə>�~)f���KU����8�[-�ЃY��� ��������$����f�W�8�p���m<_�G�[7�A��P{O.|�~��#��ik�����bʨ��Z��T���N-ՃJ��U���@�CV�-�mP����yU���$���,A�Cl���yd&�'L��=^�Z���ħ�G&.h�	4�ۍ݌{��z��0�f����*գ#	�>��c�sP��
O�s�F�����R�s�����ܡK���b��!��r1�D@�L^ɔ�7k?�#�N-��|܉��]���(ғ42�y�T".�;�"E:���3���܂yŃ�ό�Rۆ��s^�}���3T��
�uG�����_~�p0�n*�ɔ��pl�K�R���`�H �gT�����	@���*E ܇���2��{"s:��~�}V��?6�u�AKW�{@���Xv�7
AivEQ"��B��T������I�I��]'+a	�L#����U3c��Nd�|?Aw*�E_�o��F�A(]7�GY�#��]���U�:�v��.K�d�1�@G�ԥ�9~���H�G����]f�T��r�O�3���O�����%{BU��ղq.�&K	��v3c��\Rw�fH��b�e��Z0v,�l��G cP�K��N���<��:z��
�Fj�!�r�(
��;p�S��D���x����k/��fn��8���5��\��Mv�_e��sF��\SM�r�X���1j�k������*���=�N�,B>�:�5�欏��1��Ep��۠y) [��(�:�O�t X��_z�%;~+
����%�F����y��A__k�cqm#v�c�	C��!�8��}x��ܧ�����%��V����cʲ�y�/�����nGƀ@m&+��ے��7j`���QH~$"�_��UD2m��e(I����"����he/�JC�5ߙ|+��S��L%,Ĳ�	��v���H>H���|I6��|Q�Y�)DTd��ĭ}Y,#~���2�櫣�VXp���U��!%Q�L�\�pa�U�p�#*Ue���sx7���$�C�r8?M��)��X�<�J)]����������\��8ȻBվk� LM�%ߣk��h��Q�i='Q	�b���s����*Wo�R]í�j��܍q�(:�Q�	(���c}��1�*�|�&�A@����T4�i���l�����j>�o��L��|��b�����r��v���� �~}�>��yL��C��SiO"QOӛ����ţ��E`�:��_2�|���k"�+g>W4(-�A��1�%�pM�uן�X
��dC#�ϖ�&�S��0������{���5
���FSE\6pg��Y~ Vxï����Ȭ ��H!��{R�5���]G_����%%7ɯ
���S$�s����/�/ȟXw����P�x����6^R��p�#�g�<��p�fc�]�f3����4x8nW{+ X1�"	��Y-��2]��Pĩ��n�)*�f��@}��;Y"L:��kj0F(�%���Q*��}�Ñt>+L��dw��hB�.�xEH�h��e�D'�CRU$�p:�^I� ʑS�7������%C�@e�LطS3�f�Q-�ρ!��!��#C �o&�R�=������r��5k��^��?H�ȝ)�$0���o� �(���J1���N&��� �`.���H,�~����q
�K�S=��FW6F+�C`T�$t���	!`�0��@�\���$�,���:;D,&;�@,��!h���ޕb0<lO�7�s�����T����zx��{��C��z�I����%䤇1Ek�1��aw�SWm�|�S���Iv?�����
)����7Kα���و���=�
��k�#T����e(iR|_9��P�Ng�.��+:��g/-����u�;�'C���=�[����k�Ơ��S�S�'����[��K�CxB�G�TX�K���³̭�`:�V,���^��*d-Y�yD�s7����l@ �#�m4V���9�{铌�]����j�o����u7�I/��4�q�*5��b���r�k�i��L�����ܔ�WV�l�J��Ƚg�\\�'Hn��Ѫ8-�]�����5^��o������.x�*���0�zof��6�XoQ��U��f������6� [8J���9"v���lCe����A�97Ɲ�и�u���I<=��	�G��O��f��'���)�ٯb�R�SO3;���ެs��KE���oW���v��p�.�J\W��m���h�N�� 9X�71g�d@"��<\+�=(�2�}���~�|#ub+!�i��_t�������K�2�>.pu�C�L�*�w���"b�>�M=�0:��3��3��4HdU�!?x������X�G�oR�zҳ0���5Ĥ�P���#R�q��
9��������#i���l#]�� �NM���
ڦ?#j�>�	��'�= (��*�6����;�D��!�����:U�Q�ZGm���c؜JTm&h`��м1����y�69���&ȜV�a�ʨ�`@�V��{	}wD���6��.1�;W^Z���l���-�����"w p��d��4�3��P�߅e�x'���q��[�
<WAy�5x}�]oVf� �_$W�=^G�"�6C���������<O�| �\�8%������0�|�9 ����	�I��E���+�9(�
� `���i�XB�B��cb�[���HX����<�]�� J�zYr��6^��UX�ށ9�G��j�Ke)���eŊ0VA���&X�
R�I��,X�Ϭ&���iK��o���S��� $!�o�'�͠X~�͎m�����&=��P�2�ۙ̓�ݔ�t������ﭦ���{���a:����N�]�m�Գw��~�������{��i��6}����񛕎��	 ��1Rf��Sgyb*?"��]�k#6�Ɩ���m8��O�b��T�����Y�L��)���~�vu���Y�7��CByO����9420�Ϙ[��ߩ����ռG=���Ϲ��Ph��3Uz�'���̪���`(N����'��:����DJٝ�k0��ju�����RP
u�����Ԛ��|��7=zCJ�c���eOb=	�.����U��������ϡ|�7,�Ss��Ss���#�7���������kL�;B[���2՝�0V�m�\8x��\���J�E�l��i����$0HLCt,��#[�YvE�.�!f�J���]��H���m��D���ٌ�v��&���d6�P��>����Z3%(�2��ܢ���}@�q1@I	�QnW���A���6�4+����d���T[[ycJ2�z�-�W�V�� NU�jL�&Է���l���j+i�#��)Sa��_��m�N���]���7��=6-P0-�@<��a�z��3�݋�D�]t�S^?ye:�/�V�������Vt�d�ݥ�E{�����"�-�ηsqw��t�W����'��D���7�Ή��@u���Ӏ�"5.���c��Ƚb�3��lA~LI"6ۻ8���Z�:yj��N1*z���3u�Z�ҧ@��l��bB�^��˂Sy��\��q�B/�%�޷F�|���й�~l�#Mw���Sw�rLvy���4@����^�)^�}�f��1ו�V/v#�K஑,y&�g�"D���L��]��Q#����$/�B`ιE|�s�:RE,��|-m ��7�`����bPlZ`����W _��b�7���*���r����(7X��.�s��e�CA������	d~O�q|�%\���S�s3���$y��3���M���'�c��3��p�O�i��W�Qe���|�u��(j.H�曨L���+�̓����S��1��t ��,�"#�����`f��EU��7�Fʣ��{DRj�Z�,�,`n6�cx��4}�ae7��3Um�8֙�X2O9��*^ �EQ�
��r�@7U�U�E��ѐ	9�PW���N��F��Jʵ!�ې��Nq�j6�1	BĻ|�'r�̻�ر�{/������pf�3�+ߊYqƗ�^�k�C�q!"˼��2�j�aB�R�J�	���"��kh�V;��
�e#\*$��BO��s{����rp���T��. }i0³�^)LoA�[5��m���N4�5�w����A65`b�[��M1ӈ�p��PP�{nQ�Ϧb��E1���}"�G�Y�ɋ���M��p�I)N�u#�-|��=J8�g?6j�r���+ hh�Ӆbv��������md������;�C��"Y�g�uC&�O�v?@x�v=K�H�>k�_蚋�n�����m�˫��!��M��,�����A
�{؉��i6o��Y�4�VP�e�y2�vop�9��4e#˓Z�F5��B�� ��Fs�ݺ`%bꉎd��qB���JM�Z��l�O?���=i��{��EG�o_��ԏ�B}�p�q5�7�wHS�Y4g��׏�2��������-@v#t?{�2߹�8���׫Rو�]5�q)� ��ُ�]���/K�x]���>~�����j���˲�k��d���zM��G�ͷ��6le�=���^��������ʗq9����*�m��JC��U�'��5l{<!&W���fB��G=_�N�u�S��#̤7o(��E���:�f��Ÿ��ԫH6z���a�~[�����ŷn:H2�m�\���o����O��`3�VV�wͤ�����y���`�z?�O�l�w
z�c���b@��,�SeP�([�&����ú�t���%���ޞ���~Ò.�p���B�੊���ƚZ��<�w��TL6�7���tw�7f�UfR�*��u�hyWn�k����Q&�Z�1�����C����Y�Z_k��#�������tw�W�qW��3u' 3�Ҿ�"��%�E�ͬ1��L���7���KAh�{C���[�,1
�^�~9�sT��5���n9+N�O���M��;�݂���J�ШH������u&�M��ِ�f�=N3w-jeī�ߌ%X�[蔌~����q�eE5H��1�D��z��b�[��ea�an��~&eD��W�͘��/��5�6�.��b���ʛ�H�B�O�j���N�7�=��ܤlc�*wSڕ�[T�tW.�/�a�v�ҁ׎��
��f���C�׫?��IK^|6"���A��	2ʒ�������@�.DG˲dF�:�)$kop��N�g�}��y]�F�7�J��=��'��s�=k�[��#C�W�W��g���@�Ϻ�~y���T�9��1+9_\�\f�q����/ݜf0��8I/��)uh\G���@B[�h�0Qr�y{�)����7��������I��?��b�ሎ�Ard7	����N�¸��@��mk�9h�G1��t�|ZR	�5�;�/�c�>�j��Ƕ:���n ^?ˎ�bL^7�XOg���H��.��Wﱴ(�����NR��������m�^o����J[�vW���ߝunݵI:ѫhN���Ф)��!4�߶<�$2��W[��e.��8)x͓l���@�'��<�^e��}�`ݯ�����'A�rW�U�2�v������0���:�� ~�	X����ă�"IľF�=���{�gN��.&ۭ�m���.o�I��8�t��t�!3�O��&e}��Ɖ�8�����{ �%��\| >���
X���/��u���C�F�Eϯ��
Չ>J�"��/���s�	:�n_5�7X8Ֆ2�<���2jJ��t�ߺ��o,'a7�C�ß�6�/G������s�����|�+��6��I>M&�v�;�l�0$y4��:]�l�n n*�8T���W��J<�VB��!��� �+����{���iE�����GO:���!~ё!�#a˕c�0�����Ч�8=0Ȥ���[oА*^F��x��R�>US��M�]�|Ⱦ�z�1c��m*�?7�����IS^j�[l���g�yP&���4;J5I|7N��ʴ&:U��S�YmťM$#�I���b;`5N��=��Q���:[�i:hI�H��>/�\U$�.v�L�l�wO��j�r>��r+Z�'an���-�����^�hs�ΰe?J��m��Pj�n�٤R�9�0y؜c��p���܊	1�H��i��jT�vð�3�z��8��`��[xr�D-e"�။R��	�ޚ��Gsz��[ӄ3�I�Yt�ܳa��*�r���\@��ZB	:1<H�F�h�bj��'�τ9/x�*/�H}J�]cCx�� �lI0���q�Y��Q�s�E'��.C�]DVpK¡����=��T����^���'ҡ�6Gm���v���Hm�g�x�@{��9��3�>���Q(`gc�E1�!�����:�g����ge�#�
������<'�Q�^�3�qbSTF���ș�w�Bb#�͝4�>� ��2t�.�yW�T��1�8�ٿ!�B(�x0j�	�����h�z�ɄU�+;�?|��l2���5���q���M�pTvK�^��k4��D�0/��"�B���w��iS}4�7�)5�QW�0�zE�;����~�,c
�k��I��h�R�x���_�3ز޷>k���u�C��1�ۡ��?�	_�XjS}�BT,���^b/x��p����E�����o����.mN��8㕦��a��X�z �_	z�ٲ���0�EZ��'9�Y��l��#U���F�O*0�N>J�z�0q逮x���`�P+/e4�I�;,���+a�̈́�v�a����E�R/�lk��.f,���RBicJ��-��s���@s��<Z�n��M ߕ�9�(��Xp��ߙ{�A��݆`=�����_6��V���hm�@\�O���l�9�K��'�"BN�!0�۶odAlσ��r������ߎ9�R��?q��Қ0��ld�]���1(%2�����gE=���i���8��u𘳪�0$1�l�g�3��^���(=@�A��P|�C�0WX�8^��Q4���H�5��.WY0�ہ�5��;�Tv���Y�}�I����(Ջ�'B�(�'Ot���@�+
={�l��-�^�"[�Č�-���V�҇���<���w"_��D�W�3�Ȱ_�ɮ���_��)�f�Qq����}��mH�x�q%��j�N@*�~��g��1�
�C������Jֆ�<�3jEE��T���@����n�����L:��0��٨�{P�ɘ�옃��V��p{SX�M*��K�Hdn+���ֆ���9�nK�>��c�2B�锓���t�:J`,0��PS���'�HЭ3O>�%�4��wJ�|!O�E*B��Ϻ0�;��P6&��f���$Qa��Ц�_yE�|��Rˠ�#c�yw���eO�a�yx^R���(g}��eT�D�����Q�>�������F�^�@0���JC��SC
� ӱ��-�������]�x���Dp���e�l@���O㷡B/.y�7�hG�� �3��yY�j-��@S�V�K$��Tz3�Flu� �����RT�E`3�}�i5+���!a��ٙ;��.l ���Z��e���R�b@� �<}�jY$�!��@����y�v��5@,y��$�����j�40�!G�\3����ŷKQ2C��SӃ.N�
)N �cg�E|1Z�m��~6hP�X1A�ȿ�w
R� �L��`
��0����!_X�c��l�}?4;R-0i�P��
MSѨ�Rh;�-�qk��z�끯��lPUV�9�N�F̂wݷB>�g��8&��f�PBY�ۨH��y����M��vRZ~��R&��4�)>�@��$Lz�_���Ҳ�S0�o��%`5�ӂPV�>�X�����"S�ɀ�@��<2�1؊+5T�u���l2v�ӗ�B��$�d�<l��։*��^a)�$�aP�Gl@��&!�C�Cx�]���~��@��_�`��99�u1�.dvn[A=nd���B�`�qY!�$\�,]oL!d�'���������:�ϺWra�{��HU+������Z��<��VH�2^6]K{���˂;+��}{ȸNy���5�`)z�3z�69u��i���0Ȑ�+�]e_�������G�۟��.�b���h�����Q�S����ZX�b����$���]	�g�$��<0e`1����1?A��j�c�{O`
kqf4�S�������Z�J���D%��$=�w�(�	ԑ��̢Th��	�~#���[�:z�Fw�^�2�;�k������$4ddvD��*3dX�wx�CЏO�/�����E@��L*�_�]�F)�����<�e�]����Mɿ=�g�c��<nb)�&�?�e�m���ݒ�٨�&���O�[��U�2�~Q��7O�hoV����P��bʺ�d�}r�#�[(qt6�'��G�>�,�G�\y{���b�dH)6�f���[ɃՐ�e�j�L����� �/�Ί��5,	�}�z�ESSӣ������q{�Xg�0��<9tF���(ռ������P�;LT�*����%��e{�{A�UG��A���3������,$2ŉ4�5juf�����;����߬�T����^����v$lPM��w���P/V☒�K���4�f+	��=a�ņus�D����d�j¢>���Z��Ŧ�[�3^�1.�e}��ؚ������g?�����<��ؘ{MM9a#��D�����G3J ������8za*8?ן%���n�Z�2n*�Ⱦ�mb#q�����-�V��Nϖ� ���w�;�`	��(\����F��P�̜�"�ִ(j
\�]������g"�Y� ��/��&E�aNZN�m�E�!����������E���5%rf����cJ"!������úfh��]2�c��z8L������[D���;pW�y�5k��9,�˳an'��*�=Pr�r�T{�5NC����;��4�(&B#��!?����]M�u����Gn8��M�pɺ��+5Rs�O���O)���(��aC0?�"o'�]7�Y��#�/m^�A�=2*>�I�A�=���䲵���z��Iڭ�ַ�z��~��ƕ����+ϟ�V~P��Yn�"5�$�J��7\k��%�c`�'z�_i !ÿ���,�Xn�w?l�2�;��l��8A���;��/!�+^/�Ԩl�������jѴN�%%�H^�y@T4��g:�����͐_�u��0�]�2��ג^����J�ԏ�[�3׍uRS*O��V��L`�${���[��}�l#sX/B��U�#y\Ǵ�_�q�uzH�V�oh�;�1�&���{ܸ�	�h�2vS��L��L��5e43��J[T�5��yU����tnf��lrn����#EV�t}�Q.���"�ۛ%.{t\+���º�{�Ȥ�!U �q�����J�gx�H�s�!����b}���ahq���{un��%���K1�GX�!�"�h[�/M���{���w�д�x�8�BC��!�o��c2���rJ�^Z��^��,'Pt��P���^��}�u����h�[�C ���^����J���7o#e`����=w��Qh�軹~]��;���}���F�]��4�����������n���fC3�y�;?�uVrI[�N��c	�*:���T%)�1,��ߍ{P��]�>P{#ƲVA�#�M!0+ߘ�k�Ս��'��^�އ��Ḣ�G)��x4�4�=2�����0Q\�3RRK��BO,H��R(�!�[f�@��kW�W�eVN}g�d� ,���f��Tr���ڑ3�!���$P�� 1�k|N{(��m�:dT������+\���L�#G�3�d��"��y�9-.�u�s��B��3�Ւe��O&[�r��Z4܉s�kvQ�R��@dH�]k���wr��]�^<9�o�<[ߢI��oi�k��s��mL�5�487de�j4�.Y۸LR?��#��LɳϏ��;�֨\����*�y�2���k��3"�G�ޗ�׎i��B��;j����CO~��fY���<d����?_�{�>|�m������E�^W�'�)�
ƪ�H���AS�B�_}x���r6�Z�_�7�eB)i��:��o�l/I|�:n��g�r���{M�o1���c��̒��v��?p(j����:�()<���a \\�`������ݢJ��}c�՚�V���{��z_}��)�A^�$�4�,�O���#/���]|��U2�a~� ��� n��N�."ѿ�oZN���0��fڼy�q��J��2-c���O��O��\Vi�����ni��?Ҳ��Z�� J�S?U���sZ�}��ُh�ʌ�1�'�N�5sV��kM���>�8*H�8�;1A{�R�����Rr^]i�"�f����n����h��1�q�^�9B1�d�-�Y�0F��>��͆T,`<�D��'�1�^��2�Ք^H�w��7��/&�
,jf��QǸ�sN�Yk�Cާ3!��@�u3G��i����	��<��O3����Aиi��p������C�ˉ|gf_�����6`��d�Ծ�\�S���ҵ�"�I����9�c�e^�`G���$�����Xa��94/@��߿6����o�dH�D1Մ�t�ѵ�i�S�I��Y�i��<C�pRZ 
8��(�KSa���E���u��o�Vv��҆c�4�~��?%f+�)��I7���<��w������e*7���'�{L�����ƩI6������Z�HihT;"p.��x:;��dK���D*�ӽh���ԋ�^I�C�Q�k%FL����#�2ӹ���79�A㋔z`��F�c�c��d�.��Ҫ)����$Wĝ�Z�o�&f��w��R/et-b�q�[�R�7��>���,'B�ᚌ�������$X�	/ˋ ��!�9.�����m�0E���F�k��UI\s!��Ý�%}�F���W�=)�Wl�Ӎp��u~�+�3b��'�_^q��dvc ��r���۵O]�qe |�K���\>l�����h(�irn<N/\�h��u;gm�5��'�ד,Lf��6��D��������*�f���<c�@d��|�*T���buY^������*d!�E�*/3��e�����{�|¡BW���'�c�7C1���5$��1#���^�R�ˎii��?m�*�tr�՗Df�̛U᛽6�Oc�~yy,BQ6]+�xj@����xw���R�(p	�gKM�p�bV_�K��P���&��q�U��q��j
.� ��5�`��Q]?�	�.�3K,�Y�$\a��j�yw9�%2�/\�,{,��Lo7�_��lH��j����א�K�dX��{��^9���%8���<��Zb�Xh[.���1M�����I~�k�:������Qn���Y�F�iq�gˌ��}���݄��(to�w.�/,~��}q��Jt=��F&N�+a�2p��g|���ͰL�'+���tug���'�H�՞����1�I�h]h�P�� ��{Y9K�o٠����y������=��u��x��;���s�"k�h�߰��0Tqu8Q�H��p�S��$_Gt��p�^�����d(u���0'���r).
���a�ǴP�����$�@ť���\e/y��4�9���E�.K}e��9o܈S&�.�%���N��ʦv=*R<�bԣ�!�nl�0����)�%�4��,NV���iS��N�FV��aTh������m��n���"ٯdHǇGP�XKU�=�^L�1y%S�&����v`	k�)]䡳Ĝ6��~��`���>hiH=[�^��\����LAF�]�W�E�dýj��Ub���c�g���U?Z.��,��y`�ͦ��[�sҖ�K(Z��Wm�ˎ?�ҡ +m5���W�����sR����G��)p��I�$�=yyǾ��<U/z[0�-���{b�9���;� n�K�	ʠ|�p�<8ߓE�+T��#�Ԁ�,�����Ô\@ʦԚC��%��| 8�SG:_A��;���Y"�2��+�Qb�ДNV`��k�	���h�a9W��~����*7=��,�N��&H�ֽ`�H��x�D�����k�ׯ�lYͬ�Ѫ�
l9�+M��|6��u.A���KZ�0�&�M�~+��ڇ�U��
%�����%*����nl7���Ś�l�y�����P^]�W�IoM��7��y�}���R�y� w�m.JN��B$��y�ݒ����"(�ZKr��8�4n��ٕ�U��|�
�����29Gy3����|��oY��A���gn_N��-lr�������<�Agc2V=� [<���۵)��s����ޘ���%�J����O�³�{���Ls�#:p�8�e6f8�x���zw���J�?p�d�ͯ�����a��p������Bs�է ���-��+�����wa�1�O����s+z� �x�
��)�%���uԈ��Jk���K���K:y�SE��
�' _�G�A�uᴋ��%�����r�$UO�����g �Z�(>٭�h^�	�>�v��\�����-�&�H��r���Ch~+<��&��8�"������^N�\Y���o�^�Ơhc�0�v5���2FaJ�*�i��	�hu�~wZ�w�H��Ԉ)<, ���7hٺ�4���z�x9B�,hA]��F�D�Nm[�i8	��t��R�w*i�9�a���T�<z �9c4B��8��6�x�-�%��)�I���=�XZ�R�_�m�!?9ҧ����u�d�)�6�l1�~�y�*��i�e�`\�V[I-�#q�kd�� 6�1�G�ճىT�&|8N�5�����!�&L�:�;��B<rcOR2�<�Z�����?ZZE��q0w���=BՆ$$Ӻp���(��PNtz������i��`r�5IK8�Px߯C%M��Օ�S��a���BD7��M�܇>Nrox�m�#V�Wm �N6W���jS��Y�<2[���ê~�Z+��7�"ՃD��ǊR��W<�X䉧�08��m�s�$�9�o��a�0�Q�o�uJ2�C���}�AV���N*��ui{$�E����'����v��-6?078^YC��� �LR�?] T�� a�r�,D�q�s%gV� ��|ـ�6����(do[k�lz4Q�!��?<�N845ӕ|�l}�� �()Z�������9���#b������H�i�����c���To�	����5!�ѩQ��-����l�H2�/���뒪��z�!}��~a� ���[/�YdǬVW%$.�4=��h���0��J�E.��Ue��;��� ����-*��e_�o��#5����)S����;N�.����0^��;��'��#���^��\��U��hA�D��͏��T�{�1��'�1=�q���G��Ҁ4��!ǂ'��s��[!��OF��{J�M12����.�a[ٲ�=�lY�Jo���*�P��������&PU�.�b���-�8-��)�
��Ԇ�ʝ�5Y���n�	:>�w ���N����5�{�#d�0E�}{bU��[٠����=�}-�F9�F�`B���{�$*�����NI����j_9k�,�2����.�V�42��Y������� (&�;7����g[س�B�����]�kOU���&_��+��2y��sۛ4���d����Z\��\5�|b�==/��_�K/�T�8��Fg#�P���wPǽ��X;L�TD{�ԧ�@�%_���_4V�DFzp S�A�C��dY���2Q|*��Qt��+=f<���u�p}����#ۑA��<U�2��V"��CY/r1۾j����p�u���<	�5�����O�"���(�y�)�AwV�_��d$|)r�э��򳨮=zJF�tn���2�߻�՘���K�vײ����U+�@��ʣC|�~Յ�y,�r�z��'bWb�-n%0KUcHP�ڃ���e?g��7�bXq����.mӮh��6���E�uC)r�c����`�'���s�&���s<��ⷼ�^�_p�Юs�����3 ��)�6
d!uA���zG`�ʡg!�Y�]�(�x&�Ƙs(;m���t���\��ד�R3�.'���)Aq^�Y�6\�L��k�6���+G������~I�@�K>��* 3%"<f'�wг�O�s� <6C��r���gZ�$F}q�[�j3��{��z-�/�k�m��TL�����-K�YM��]��J�pt�B�^��~<�rQ6�P��՝�Aѡ� �[�cmc� Z���J ���ɵ=k��:#� �ݠ}�ט�
���"��F������q������V,2�ge�%�nn��aB*�A�nq%��3*�7hy�@�m��Wܜ2�-6�K=5�nC�U0�0��ߩ� �?���J���
}ۚ�t�l��a1`%PZf@���a�wn�Fs|����檃t��<���K�$�釧4�4^���mP8R�#�%��?�/6�Б��J��`�~���	�����魯<u՘��`븰��t�	?���[2��<S���,�?T�f�����x���0[Y޾v�B0��H�k�|X���h�7�Ω����n�N�g��Un	�#�X�ɶ=�#�L1�	�}��x�Ջ�~��Q��_5��|�jXn���4O��������(�=�
 �1�,����#[�C�ۄ���eQ��=���:�W�+"p��@��z���œS��瓕���`�xT�Xj���s: xJ'�����?Z��\��IR���߾�M���_�c/ZEF�j�OX��5��?ue���]���N����y*�]�3jL��k����C
�k������VngB�7��d���{��M1����6��y�6�|nZΈ�J>�>2���=��y�g����M;�ܨ<�xe?P��^T��O �H��X'+�$Q+ �	�L����ض���\�\?}m�D.V&��p��L散�^��n8U�cљ���W��`)���\^��_u>���g)���w0��-�ʰ�����2�3΀!��ZZ��6�!��h�P�Q���Y`c-!�|�0��q���G��Hڔ�AK-����m����<zH��&;Q�3m�_��}t�:W��5�S�l��aI�:iS��:ec:�_��-\�ZQ�ؗ�\���K�u���a_�Ԯ�)6TB�����Xh�}��ǯ�+���|w�1Ҝ���`���@}�\Zp�23^^�ݳ�௭��G���W���i��=�k��K�\������A�����?����~wt$��'%ϱE8����}�J�@O���a�7���9���\���^�̯���g�xd��alD��1FD��	tg��n%,\C�g!���h=����$�[܅�lTj�W�������i�qؖ&dL�$
h�g�i}3��j�a (�g'�F����m��3��2m� �o
���/���&0�[f���:��7&����\R$�-�����,nv8;�3��{9�q\ʫ�`I����.W�
!�����7�ɳ����'�)gC�OS�=�Î��q���a#�4F�ί\�01���ά��Z@���JMΪ�%ۮ���'K�ŚϺXG���k4�I$g��^F�Id�2L���+}b�k7�{O�/\�*��EI� �؎j���c+� �\��#t%����R��q�!�۲.�|���@���7�1�D��9�Bڣ*������E�	���	G6�,�r���؛�q�1邼&�Z@���Y��<,�  FI���MU.����H�m'i˳)�\*`��t����E5z�|���0^tۺ�t�A�>^z�<�y�X�:[iX�]y��o�3����>l����x_����C �D\��ݝN���;go=?�]2�索|\JxZً���*B��Q���gsNeO0�Bx� >��=9��H�5���n�6��Õe���6��JC%�G�=�-�0�C>��%\B�.���8%!�߾�w,�}��Tg��p���d���J�F8������4O{9}���)�,�0����:&��O�/w_�x͑F{1�1�$y��Rڵ��#V�k�|#��_�_��|׿�,�ҡ�K �n�zjs{&��=���L�F|��DG#+�l�W�<$[l;���hș{�I	F���'���UH��)2�� V6���8/j\7R���,�b��o���v#�\����TS8����(�p�`'���lg[|�K�8��p����Ω��g�꒠�ˆ�m�g�I��Mw���.\�Џ����-��)(}�2���j�z�mY9-�b�$�C�51?�bo>�������//���GhBE^�~�$�A�����n� ��vj�B�U�GN�>
��W1 ��I=�s�o�5M���_��^��������	4��W�l�7Wɜ�/7)��k�;���4�t�K��S2����3lNO����3�N=��ق�0�]�N����Fs�ָ�P�L�h���L�י�X0��6��\ۘv������O���$������i~9�RK]g��Wu�l�G���ݳ��*�� Ɉ�Vĭ�9xɺ֦��T�O$T}+�A��#`������h�4?��"��m�"v���d���]�q�Ӊ����),�� �O��Z��{_�s~�m!��G�{���\��� �R�s����Ϗ�%P�Ҵ�|ȗ����.�D�'���[��Tf!��+� Jҿl��ܣ�h�Py�W�z&i�������?j2$�&�6��䢐�$���9s:�Q�k���J새U�2�����Y��S�D�����n��2���*�_`�*<䘵,�=n�S�r��߮��<$�,2�$!���:@�Ԝg�Ѧ�r�O	���|�S�q���]2b�k߿Wyҫ�(L��%��Ļ8�U"NȾDǹ3ѱ��h2��'9��.��1�3�w��v�~�q�����!��ѣ�񫱋;�� �۰�@�
]��t8&5z熚(�����vCkm�I9���v�Y,�r�dN���Y�&�.��D�͙�q]�h���Lx�Ts�.mFe�8�E@�ђ�}���|^v�f����"������w��v���D��~�	sAݧ�Ñٗ��_��&�C�H�
����G�����(�g+
�}5�)g��-Y̓,�>�ާ��؎O�]�s%�n����,^�u��Z֙�V����~ri����
%����_�a��R�.	ee�J�澥�ʍ�������%�]��f�SH/�].1{+�������i�@��J`����IC	�S�i� �Zn�xA:��(,9��Vħ�	G��pe��(,�9T�$ �{|q8V���Z�!0-���E�_��^;=?T�}B�ķ8xc>'L���!}��4r�(>g�&��������'����"C��ړ�e��|s�F�7������G�EU� �٥:��CzW���;�m���r�u���!���(^���T��φ�x��ߍ�o}a�� ��j~+<���P�Y�ؘ6�{z;�ό�a&�H%Rm�/�y�ϙ����#��=�
 H�ǭ�@L��۫�zM���Uc%����ƃyr��*Q�!c�y_C;�uǿ��?���D׍2�΀`u��\� 㬃��z?N�S�5k����{"�̇̉h��/��f�J�ϧ���#ż�c��ϋ%_��xu'��9�in�j<�H`�Eh������N<O�v��k�֭���$�d��I�i�*����Ti��"t%�Zwm�V�d�U�� b�&��1�@3���:c^!� 2�C��8��/@s�p��8g���yO��I����>�Z�!@�R�����8
��;OZ�U�lf.��b�Nƽ{p�ý4	K���:�P'#PՕg��u���'h��Z,Ns��o	�Nkga���8�9$>���I]΀�Fү/f�t�Z��=��'����,b+�U�4y����h8����M�E������3�4h�o�%w�42�fOeK���7�q������d��a�I��h�+��Wtz�\���:��'���� n2�Q���@��Rf�r��h�c<v��J�9�2 =����Yu�Z�ߝ�_��'� Ԣ,Ϧ"4��H[�Te�2m�6�fw%�`�' ���@W?�o���]�M�H���;DC�e����e��&J��Xx���o ���<�����=j��Y�?4p���R��xcm��^r<O���翼�Ѕ����.���z��']"31�>&��z�z3�(h�z6�DJ�����@(������ؖb&?.4��h��p���k���qgj~]1����u���B��nHf(q��-��
p�����h,��QW���¾w�Ei������OV�L �B��=���0�2�vTI3}�I�18/�(q�����(�B��xY/�S��>���ZDS�C������EZe�8S�W���ӻ[&A^������uD����_�ZEGA�?\Y�<�>'�Q�(�n��8,HM�l5�N�h(���S��x�¯��@�k�M�M��ɍ\���=>�O�=����t��_:%�����P���S[��.��jײ��?��m���P��N��)C������y�|�)ĩ�j�)�ɉ ��K����U�Q���O�E�^e��i7�
#'7ɫ���="���� ,�8�퀾�:#E�ݟI���Hӏ�y�x#&�QW�;��M��U{��9Jm39�߇�$��C&6ؤw�j�4o�ke�|�c.�a�1D�	1�>����m=ti�N��?���@iV����ʩ�"a7:���U�P��7�K�/2+��#°�s<����.7Q���1^�����ފ�GY�}w�dX�[���weS4�[� ����U����Q�	p Q5��.���� ��I�'�5�G��l��ʺ��2H�╻D�u/�K��P-.
q�le��"Wl�6"�!8j��ѣC#�zC��>�1ڀ��"�5��=Խ�v���Y�C�1t3�x��������rv5*��!(]�O�|md�
�A3��h��}�t���+�J�,H=g�o�Y�����\Ɩ��&Y@�X��[Z<6���M�֨@I��o�p?P�3)!����a�C�8��^���8��7ԗ�"��?�%0�;�cߑ-�A��ŧ��>M&����n
�(�Jѩ`GzCkU�[@Μ�HJ@$#y�i1����|e����-^ެ"��_\Z�6Uzol��Q�&�T�<��_�X��u�a�5ОC��}�; /���}t��2[�����C ��T�Y��UG̳��
k��fM�-�]�@�V��lP�A��Z\<̠&֌���#��o��>�������̦H�X^);p����B^T�E�;�%�BnM���MFj��J�RD(����ڔ��4%���!���Ȩ���xy�j�8t:p-�;YU��8!S�^tCT��{l�mM/;��6���Q�)4�86����?i:�tT@sʀ:�t���zآA���� XRc���,�0FjB�|�.A~���=�]D��b-��}�:�D��뵦��_u����&���b�N��J�+1g��!3�b���<O1b��p:�����@|�K��3LW�u��*G���צ���;�$�zʹ0徃7�v{�8���7����B-�{2���ȣ�����i�Έ=�x�M�����n� �վ����tJ�*[������&�;乚$�Q����'��k/�hb�	���H����c�ٔAxv��� �Ϭ$�K��Tq�e	��M$����6��f�JQ]D<�؉�������]a��V�]n|ٵR�;�~L�a��JL����uN5�A|/�*@�r�K`wVe��;����P���o�n��G�P�i�U%w3H�w�4�����d�(�A��k�\��K�}>�`���A��^e�i���]�G�ѼB��.�w�,�������U����v��$��~��-�K# ���obv����SϢ�?ţ	�(�\a�)ʢtp��y�2Se��4�Z!b �T��0����x::_�IU�+Tk���2N��P�A�"�B��i��N;��1Z(b�m�~�� /����]��)VEJ�^W�p�P~����֘Ԉ� S,;[1�~&?��L�=���clN�w)�I޷>&=u�'�Z����x6���z�����TS�SDo�~�]�������4v;vw���͚P_Sn�����Ԟ��vۻ�9]<�nq3Z m��A���2~�p�9z�p�0º��wm ؑ��A�$����&ѐ�������W)���{�AAI7�3�}��am��7��м\fm�r8T.z�{`?c���er������	�3��}������v�"ӴO�A���H�ͪ`��ւO:�T�*#�Cq�-��:���/5�u���������Mܵ& �Ｕ�e8z)��\7��D�=���6N�G	�V���W���4��$`7���B4��o�h��t}�y �p�0��C��4����gn:c���3Cn��O�}1'�D��SW���+m47��w�0�`K��=|5�0e�����s�]�$=�BV'C\�%�42'�� �z $��*cr	��{8�������]�$�5A��w�eΎ�l��{���2���A���+$t�������� )<Z�*|�8��YK�o��f�8��pt�����~����Kx��m���Yu�Vbϋ��kZ�k!��1.8��aÃ/���[Fr� � �B�v���
�һIے��"��@?��;��MmkA�9�W�ߒ�W2;�{�,%��s��j��~��{��1Y���M�F^�q��e65FT4y����L��Z$� aqӭ�C�[��yW����uwT�Z0T��gY�G? X��2�����,|�UCo|e��H�t��|7D���P��xt/���M&�<	�ӕK��⨙
��+�N{]�ᩊ=g�=@��1�|��v��.v��͌
S4�1�s�W$<��̝����p��4�83|p����s��déoL5#3��sH7�M�e��sլ��n��*M��7���� �Һ���� '�,�q�Km�7��@0�}h�
�O`�Y��pj���ֻ���{}��U9�M!����.����#�:�I<L���6S��l(�:���{g��|�`����׼(x�a���I��&@o����Db^���h���_���?�K��	"�{}L�_��|HmADS7'����2��C�k��[��0���^H��ts�=B���+,(����+�4܁�<�S�%า�4���:Һ��oXJ��PuFP3`�����ǧ<+6l�fA!V�ǦI\�/�@�af:N)sj��.3R�~�\�0h#��ǰ��b��2�ʭFL���^ƨLr�D�}+S݄$t��0W8��bs�D���z��d؄L88�" �^���f�P�+�G��.��5�V�j��C$���%W�P
��[��
�=x�e�^_���a�d�G�<(\A��!2�uã�,tC���WܟE|ƾZ�8�ˁq���� Qo��\��(����oD��F��^����ލ�����@�>OQ�>IaG�d7W�ۈ�������.k��֯��y����,���ff�{�m�QF@�$x�_� <6�Kl�p���� q��⪤H����A�>��Ø����B��`��!hЅwɯe�>��Apf�,xhi�Nd�N�)B��2�+e���w�8�
�>�y���:0���F)Th'U�E�?&Ƃ�O���a�p�G����m��(����*��M_ߨ���O�8�[W����g�W�滤�4ύ\?��d�5!��b!�+��b�E�m4h{��Ix�=��Yny�;WL�z�/c͘�"���E�^���uk��}��\ƹ�C ��Xe�L?������)u* M?��;;�/����H7�KA�r�Y�� ��8�!?�QF�"��C+��{,�	Q������n���T̳r��w �o]��-S=]1�m8f�Z�πV��Sl�|�(��	~Wk _���� S� YL��q��ǧt�w�H�O8&=�Ϟ�;/�q�m�iblZ�%�ѓ� ��GER,۝�X��l�n��L��)\��W-O_ي1c�I
Q/J�O�Q��A�W[|�c�;͐��ަ4��C�.bʸp�@�զ" ��Q�ϖ7�Uom�e���\�1���
{��eC���D��ti�h	�*� ��A��\��{���Os�*ۍKy|�YkD�#�)��@�j����(��U�1�I�R�c��W��Rs�R@g�j�0�}ӟ�|�\�e�$�a��[�����s��W���a��q#��_i25�T˗[w.3U���p��X����0tX3��ig���F�P��@g�x�q��KQ1�"�`���v(�;� ��N�ff��� ����$Ǣ�TE�]��G�*�BY�O�1=��g��W�%�{+����ހ�h{���z@$U��+�R���oE`ß���G�&р�Q�PÎ�`U���%�<q	W{����mZ�9�L�D�V���.B�J8n���� �U�W%�Sz ���7��2^cacQ��*�M����ٷ���S=M�o�%����A؂����O�uxY�mkn`���#x|p� H�V�7G_��銼�9I�T�H�)���D�I���f�d̟+�ɬ��i���&�Z����P�7r��Vy��D@��pC�n!�J}۹�A��?Ɛ�j�B9�呈�d�	tF^�NTܛ�S""22S��W�Sel#�	��
wIG4�?������L�a$����:W�X����F��W��@�>���zr�"�W7����9!<��P�q�N*���"2�q"+-�=ь�\��+��~�Y
��&�����^��"�&/��22�r���1�/�h}��F�v��j���<]Q�2����2[oI��B�*�.%�o�{��9Ǧ W�S��ˈZ	�n�k�sԕ�}�@<R=_�������􋋐�Y�
`��D2>�,�5(���� �y��Jv�#��D���e���Ƽt'�H9�5�/4��ա���Q��w�!b�����r	�s�w\ê�D�Pfjm`&�q*�|�չ��*��]����j���l�?��FP������B�L{�9��7�_��D���G�2tl�Y�m�MIq�O��=0�BΧ�"���T�Z�r�0~{�E��zs�ک�14��M�$��@o�a��ɿ�W��+��Fs��KҢ�������1�IQ���$B_KC�9�<©��d�J�:�Q�+�eȜ�ET걺HL�T�(G�n��^����%���\����OB��7����*�� � �aa�J��X�汭���5srnGo�n�KGS�n��F��l�5������7��zvUgyY� V��@��6��-s�X�]x�}:p��"�b��_B��p�ʇ=P�tM���t�)� �	&��V��?k�c1��{2u���&$�B���_���L2��)�ɪ?��G����f�!���@Zߐe�]�d�,xy#�+�Y�wU�L��!�}��B#�itgf+L=��,��5��z0x`��Im��fD`��������7�>�։6!9��S>ߞ��s���d=�������r}�~��%F�#�����9�*�����S;�o��C�5�Phw؁���i��ŋhsnnqT[�e(3������J�6պG�ꠙ�*�҅�Q[�*T	,~Y�>wgʜO`oy��<g�2)��I]�GNR:���,q*�Ge����:{��3�1�访�N��Ʋ�p�-"k]��˶��87���'�K�aF��S"�7w�ߧX��{6<s�e7��o�yjpԥWn���*q�m����`x�Z�W @g��Uf���j�KZ�2�^^	��,yH�6�0�Hs	mY;������h�[�*Ν�	©��h��įg����ǭ̂�:��%����_V/������G�'�U0��Zo��*2W�h�ӱ��k��|�����Y�͋`�gYʐ�K�Obt�\L�d`7�/*�E�m��:0Z��Cn���l}�������ym��qC���K�XV�6����O<=���*�6�)(�k7i�s=��h#�Oug!��q<�;X� Ǎ�7���/���z�-ԃ��R�d�Q� !�Rx?�q��K�<b�P����3��$Á�r\��`޽(�F2.��99S%H�V�B2�p���9ν����{a��짡n�ǐ����r�Ep��k\�@�g:"-Bb���"��;Сt�������O[DFG��mLZ�۴*�k��:.kN{rd���=��P��'X����^(	���fT�A��J�J�X3 KY�A�Zp���Lk�M�C�A��Ԟ�{�g�xR��
�idC�/A��q��u��Vu8���t����養��_0�J�x��:�dX���zI﹞�i���ܣ�:8��^ŽC@,4�x6�4�t]�����|"	�T���IƖ�.�u��FZ�j4����$R=x�ހ]oD-r�Hՠ��c̮��vzL��/VЕ��m׎��!��n*�'`�%H��lv˷�T��lܪ��~�l@���`�������s���{�����h���w�]��k�nl�˜��������f�p0�s:B�q�nN���¥/ >&�58�G�sP+��an���X	#���Ƌ=0�����Ǎc�B�����B�.�8�k�*Jjf��/�*PDב� A�h�I�%�hRvm�����z��l�K�pz��$�V�W��c`=d2�
^��r�Lx5ȅ�k7�o��};F׮��p��CB-���S|��Ǒ���$�>�ڈ#;b���|~��Փ&�qu��͎IX
&�^�.��5��c�XY��`����}�g��W�64�J��� MG�n�Eӹ���ؖRU�j<�?cgОP�-yFN�<7�,�ĳ��װ��i�t1���VӲ/���G���z)1���mن�m����JJpx�Cֺp��ً��5u�QU�r��s��z�L�cL2~3?������Z��
��y��������[C��k?�<7�����>����L�$�>p��#�:a�`RΞv {�4��g�"�?�������ӌ������:�Z9~�iOxJ]����Ôʹ>��t��L���F����p�?�����a�{I(A dJ_k������5P�I�I�6��ARj��k�??�h%c�3��#1^E��O����|=@��y�m�7��}���^���+n�
�A�� �t�?:�� ��gQU��t����*��O�K�/���J��b&lzx�d�I���Xu/Oo3�ј��6��%8ڭ�	��ѱ��a��ۡ(��;�z@���F�B������`sV��}����r��#v������>��͆0V*M��؍�^WP�Q� �p
[*7뜷/&������gu��.d*��"h`��<Q�|�غp6y��E�U��8;��+0Q�NJ\��h��g�j<����#���6;C�4su7|��@��4Z��c�7@B�K	:���Oj�>����d����T��3��}yK�H�'�.ʫHx	9M77iGl4vr�H,;��J(����_���-æػzn�εS�C-Y��hM��uم�1������}R��Y��}���O�L��Y���[�:��ŽL��=�:��MZ�gW3S�Cu騁�p�ۥPl9]�d�u�F���f��Q,�A���^_�wH��l�xٰF�R�t��}t�μ����A�	MqO�@�-���ͮ޽>z����&=��&?<��.]Z�)׫�9��X&��ۋ.����@�f��[��'�;h�pzgw�E�B"3 ��`],�n����Zmt�Md�U�֞nb������
��W�f1�'i��қ�(/�3�|�1pk	'�A��}}�L��H+!M�HU"�'y�@kъ�(��@e<�I��ioI�k��e4>b�7A�3�Z߱H߇��C�y>��x ��̎�y�#so��R��ۥnE�r80�������=��J�Ja��u
@�Ah9ja"^�ɄJZP���/�� V��R���n��-EkP�z�N�Vw�j����n�F�#��#�'�O1�����6�y!�b$�)�F���3�^�A��'Zl�4��9��ݏ܅�.N���M{�[r� �'k��d�Cz�c���Y$��i�E@�x���t�h����VK�Po�274��������F|�E�u$��^�	G6��~�S®dK���ۧ�s4m��p�b��7�2~������X⹲�>�R/7B��\� f��rR��T���"��T�P�
#=��k�b��E<��kXlɟ�Gy1��H8C�!X���(t�G*�8���5����!�@
�+yDƵQKL������c��m�k��CLE7�]����&�Nć�S���Ə�*��V�A�-�/7v�~W��R�%�	g�Ҁ��/F�����J�}O{�?:3�ѳ0�C5vܑ��"F��l�+����1������9�<�&O��Nٵr�ϝ/�PڳŹ��J{��D�b����戌��|I���T۫�g������:N����'O�6(" EN*�V��Z�
=�zB8���1��5�ԭ�M�[�D���ү:�SRH~k1�)==�3�td}f�@S
��c�m8�F��<ڍ�a�R�e��m���b;�IV�v���1������Ņ�N�ɓ�F�����7!��V�Z�p֬�+ ��r5u����DnGb��V\�ٝB�Ei�y q��j���a���ƙjs��/��7 P�[9Y낾M}���1�����\�Ŝ[8�����&���zH��雝a���ؒ�I�}xo8���I�0K6O�=���+��hq5�K�&I���M|���HI(�QS������1 2�r��d��JG�c�qI�xX� ��QD�*�g\��e�g�+x�s1���̓�z?ս-=9�hײ�e1ֶ�c���Ă5!L��*�� -_��U��/Er�=D�2�cE{�
P�`��Z��b��d���{ #�p�Z^ӱ04�ӆ���	
#�J�;���p��O@sAK�:���L�RGf�0r�O�����&'D�9,�aHb�?�ɪ�x�ao��������gf�V��:r�[N P���U�?'�1t�ȭb�3��b�{N�rNo�"�˟��x2ɬ �|�8w79��#���{���P)�)��P*���d[Ļӽ��M�A��7�)r�OpGa�sp0�� �
D��f�)F4����0-���+]�q�%$�&��u��(*����>��t�H�JI���xr�J�GW=����M��ge͟�k��,�e��k�L2	Uz�s�j~�vM�`4�X��@W$���ЩΉR�l�}����*��B2W%	�D{�~��x�Bdݛ.Ly��d�m�Gu����#�N����yuO��p���&ȝ�A&EI���`�"i�(4�t�rcU쒲&G�QA�jdhF�ﬁOq���gպj��������o��g7Rc�+�B9^\ƽ��dSe���ݜܤ�gʍ%E I��iM��j�Ly?)��']{fX�+�k��wu�+SA��<���� ��F3__��Z=nLT���R+g�'��Y�w�L�g��z_��_$�[�H�8fͧg���_;^!ǰؔW!��`�$�~W}�%�3��� (+��u��KK�#�����S�	Z��!4���h��q��ݤ�O6A6C5��� ��б6B�P]�)�lܨD��rQg ]�t�*��Z6>�5*3VT���G�]A�������GZ�Q�a�%��S��/��-�Am�ղ��7�k쵬�HmEsGK������Jg�^E��O�BIp%��"�"���Y���%�v�&?�̛j�Sd���F��)rܓ����S�(�v�[p���,�v�"��e��;R8�y�ujO�rXg�ڢҁ����܅	Rc��9 ��%��
0�.�u����]WY����� EӜ4ߔ��N��1�f~�mP!�¯x�L^�?�	I8x�B٥?F�0M�S-������.-0�U,>��$>�0��״K�s�QP6�d5�)�(����7��1l�	�������H<�8����
�%��Q����`���;�b��f�� @~~/	��a�j�#���7�F�LW�"�{��M���I�-�6�F�D�j���*]�&��jL ��\|����pLSS�$��z��L���N?zO�d�����]��7l�t���
(�&4��l�Ä��@�߫�&[�1��h�K��o�6���	{,إm���ă��u�LzEf{Mn*Ct���QS��(7q]�1]�U{X��B���F�� /��5���
ŇpoE7	�,S�};)��~�[���Cl��8�%��g�&�{7���U�
2�B�����­�鍉����M�8�=����!]�B�bq0�]TH�T�d�"Du��1�Ý.�XH���A X,�'Q7]"+��czgh�������E�H��n�I,7��5��������
y�(������}��Y�ֆ�wU�j����焺�w!�:����`┲�YWp�JHl�q�+�n�jș�-T ����2O(Q܋�,Jj�m)�s�%h�إq���Q[w&:a��KWfX�ٸ[�	hD�E�о&��ã�ǅD$�X����-���6(��-���Ѐg}��8,��E���谪8S�]�)N��o�.j.����; _P��sҗ1�2���"��N��R�~_ ^g���Mf��)��>���D��+�6���h�?���6���+u^�����g4`��7Y�
� ��)5�]{߮�����ThM��� !���UX�#���5հ������q����Uui�������z�8�tP���R�0-'��x��g";}��Y�1�վ:=e��%�n9akp�tլ�Mا�d�[y���?���L���`)�@��(��ߺ uS��_ğ����z袳;IhP>�1��s�=������դ�y���(X��zZ�_T�߰y/�X	!���
�,�-���� &'���J؛YdH�
��N_<�<����1�=,qU���k5گ_)������ۆ���<J4�[�����2��O�?��Wyݏ��9Tg���L-{Ý�!��46�^�������r�R ˞��z�6ݰ�2�j��t��0�`��7k��ot}R�"�z���������U�2U�C�[	�����Q������UF�9_��ᙪx3f����BV����7��5g1���:�.���#�R��4�r�~@N� Tq&��$_��R�z�운���E��}�q��կ�>])�SJ�eV��I6��&N�cu�'$�E���'T���e#W̤#����|��th:���i(�s�۲�x�0v��Ξ�zJԪU㋼���VS�������8C��ﶂ�I��1��N���Bn"�ԃ�+�>��ðJM�����T��to�)S��U�����4��1�CDy� õ��б*܄F�(��<��&n��U��f�a��h��L�9��Y]?�����n"t+��8W�C��(�9�%�&�7�|�G gE&f ��X|�<<xjLl"o�ݭ:���LG�Q;H��)%�Xޖ�/:}���6���i+M_+K�H� w#T��%��_S���O�J>���`��+P��N9�P���O�и�ב��5��1.��Y!��@f�j@vveV'���'�Vٵ�������]�
J����eX$d�W�~y�v�7Ln���W��Ga7�|�{QH��҃Lò�C�Q�ȏ�LѠ���>rOU&��m���d*?�<��\s��#vK�?���H֞Հ�GF�}�Ϳ{��h��f�#[�#>B����O|�[}$�%*/�-��Ҷ�ƞ�̇�r�k�¸�}��$O��eY&��]n�{�H����]-�5�0�r��B��aԇ.cB5V�����Ӗ�a��q�:�����$Y�v�lP�Up?�!mO���t�|�H��aMJ������4u�G^%ь(�'��|!v-�4�m��mI�F^���D|�#�����-���:ל�~�1�UP(	/:,sd'�v�[R��-3?X�9N�#0Ɨ�VF/k$fK�HD�n3�l���ċ(�m�ޒ痏��|m"	�^{���\��!wq�9}��/��_���K��9�
�9; p$pl���#���T��ÖVa����1�$��_,A��*��54��up3�@��>���=Ǐ���Z6��$�|h�8}�? �(�Ȭƻz���o"C��y��O����&��sp�e�,���1�Κ	��,�51�v��LL��f����llQ6����Z��9p*�]��"�T�*��:u,�������������1h�"S��z�ڝ���O�ō$��ve�h�&�8�uV ��h����8�rX�L(NW���_���׼�}I=�)戛2`��ֆ�ZO�j�2Ȳ�^\-��͚zaua������G�}�9�*��t�u�]�NnS�r�K����&,UL��*������4O�m����X����xſ{�/G��	4��z���D�=ZR��)t|��X0ɋ��m M��Ӏi�IK�B u񤼧��!��3O�B��YC/Qg�YNDi�W6>���E�y/L*j8�(r'U��%c%�o�>z��\�nK1���%����cl5���x�>2�3
����h?�(n ?�ES�ɰ�+��O׋����\����ŋ�!�mt����b6P���uŘjư�� ���C%|������brR)=�7�Ҷ�L�-�KD�,JT���DN6��õ��s�3��M�	��6�лv�ep��#Vm���L�Q���5>KJJ�#�&�Ry삒0�/ƶB��w'��x��r�|e}Ug�Lkã6���׳�����N6t}�ACN P,VJR��})%� �]+/:d*�!7ߘ�
�NEB�o���	=Z���Q�0�uS3ɺK����q,��^��
�T��#z���R
� [zAB�p}��˘���:���ѧ�R�'
L�$�-��%��Fbı��^S%��Ҹ��%�o�7(���U����ѳ�O���P������sm�f��K�����c�&���@�d��3�;e��{����s��U�M*&�6r@��ȼ�J6�;¦�Kf����6��,j�q�^��ڌ�jm���	zkz*MFa	s��l3k�"ɉS�
�l~�7�庩�k�>H#`�Gw�L�BjRTⱅ�G�Uď�]Y2��2���Rq��HU�7Jn�|5��4$���*)�(�}� ��ʺm;���� ��d�-QY�۱ a���:��iF�;�E��3���V�9�g�y%�%��aN� ���f��3�
ӭ����M�
���K��Q�_Jzi�ךYySU�?w�q\��� |�ۿ�B�˰�n��N/�h��4��_��j�~���s�;��zJ�i��}@�{��O����(Œ��jP�]�*�4������C�� �'��Qw%�t6x��_�m2�f�t����KuGwn<\�O αl�%Ы"��q�b~�o�Qŷ1��(�?�]���\X�3�*��ܤƣg��W���6`�;�@IBF1A�C�E�({z���AH�o ��L�tD�/O��yg<z�� �;�]���}��.!�zE?^���Wu>��"D��ZV7�S��ғ+�#��[JB���d8���Ш����p�_r�Z\���?X�	׺(�;*[�v���P}�U�l(P`�BW�Xʽ�H�8n��B%�u��}����`"���b�zuy*ju>w�C��{��l"-��G�ػܹ�[����Ac8��&6Y��X��9	!���x�����#-A�A�l��F)"˲�����S���k�"��j`�.��m7�+0������PA���%<g'Č_����!uyL��9#拴��h�d8CC�v@N��rU^�I�{�
A�$�v�V�Qn�E��Y�͝EE�-��.]�S��Gҿ𨣿n�y��D:vJ9-��T,�$g���H �<�ݮ�t�Y�!1����$'dm�h_]8N��O_����S�br�hv�Z~#' �$w�1�Ff2+�����wKg�8��RN�Fb���լdʦ'�:��(r�X�c`���"�=��6a�����pQs�}7N�C73�c�Ӟ��Ølf쉅��D�Wuopj�a�[�˓6����4%^�[�_Q���mc��u��m8�@�oD��[ź���D)��T���+�9��'`�6��W������Й��G��B�I��8�j�p��W���l�"��N�3��,*I�pf(�48�(8X��ӳi��t�M�"�;�m?��@�"��H7=���>G�j�%)�B�u�C���'P��^:?���,�k�Y�D�=0�CZN2.�o�4'��Y4V��4�(�#)��_��Re3 ���<4n���b&�����]$s��|����0	~k]��e��>o2.2�2^�����S�����/)T�$�� ݼ��A@&6r�/��r���Q�6U�9'�d �a5���Y��/X$;�Bqm�hi`��݀J���\�JD�+-��(cM�'Y3{$�"�C�)�������B5Ox=U.����Ѳ�%�N�ǫ\[�4���z�nƨ�s���tm}�'�-�CP5�[�v���I���;f�O������o�	YA"���I�ܸ�G\����
g��[Ӓ�z�$-�%��T}R~��7#eǂ�>��R�D��
�3�Y�9]Ñ�T=����0�[�ʠo�rc��"qlt�X�[G5�v�i8�T���ϓ\�%����W�]ϲo�if
&t�>{����Q��Z
(f�
�*�s�+Z�K����O�6y�]C�	/U~&���7�k�W
��;��i�	mf��{._CX�o��~f@���F�,*�׭��,��ݰF߼(�������F����i�e���O~��!�ԌMR㜡Of�,m|��GP2���ҕ9�n'|�;r!m����bW)���r�S���Zm�7�	�*u�	0��	�?�^�Hv�Y�r�=��zd�m�z(�m�~�䫣�<{2UDE�B<&OO�rT#d%�]���JA�7�=��ox�4��7��A��R�]�������w"�⥞˴�Ԧ��w���)�] ����3~�6Kr��f�(��]n�%�F�����'�5#�
�0��鼏��g�&�����b��"a���#�P�I�79�vI犏"0܁I�1��O"{�����:`ҳ���f>���z!!��7������S7&���֔6^��6˙I� ����E��$��������>=�� �t�4����&�=�VY��H����I}���e2��I>h�c�N,�s��/�CP�<�^�m:(rr�6
�<(��@�\��s5�$��U���a�b�V��$��5]̲�30٦䙚F�qi���`N4` ����T�Yk����I�Ȼ*�V��?��5j�_1mV��k�s������i�ꣅ`���	/�|>7������#��X���7�?�����T�-�8:���P8b�᧩����$��	$-�-,=2�V��qx*�1E��* l5�-�09��Q�v��i�|��`ц���.�F��@Q(��")�0���}��-�����ϐ,��͂�H)��3�K�őت���T�x��c����[Z��qA�O��c�%L��,	Y*�f9�/!���M�c�(|���4�w�8Y{4"N�|
�{V��Õ�X���ͧ�AEjZ|�6���z�P����ѓ���Ju��mP`1��~�����f5��r/csM5��5i#�3P��2�Sx�����J���L���7�뢦o��I�lT�$FH�W��T��H���ήX٣,7z[�������M?��!��=}?��uc2rI�|o�϶L�4�v���(\�#��`�Y�D�?x�e�҉|�n5:T(i���,��H[�:�	R�;�jU��)��u�������`r\��8Ch 8���WP����+Ch"��U1��a��$t��e���Q������ʪU�q��?P�ڇ[����� י�����x�)�.*^�h@�C	�Ip&�cI��f�b��mT�K���هj������@��%.�Wn���C�w�bSH��}�Y�2�F�G��v�5��T�M�R6� MC��ywpP,9�օ*��j?��&:�	�;�Ź���qlxy�^{��CF���M��z��_\x�����������7i���w��D��S�p��pᓚK�/���w��	��a�����Z>�2��;KW>�~R�O�ص�v�
� �
:�e'y��1�Um^��!�����w�yz��ⱬSb$�Cj�a.Q�紀�ie�+uNW����16�� ���n
�Һ;�r� ��[��Ɉ��_���?���[v�]�.�Z�S������y�UԵ=<����w��Z��������v$�Lk�K�n��X�yIR�8�4��P�#���U�ƻ?~B���δ8��d���׌j}����u(��8�ȁ���
��ɬe��������'��~��.��Y�ʻ����5��$�>��ޟ�7��auۀoR�XW�c�F��~n�����&�<�PJ�@�y,�{���{q<�\릙�+���^���5��w9�-���;��WB��}o%M���^kM�g�$6r����f�.��|$5�Z�E������Nv�_������Y�c{8�f�;���?Ч��hd~U����Rb��U׸��p�
2H,%��W�����5�VEX�D�[��iV	�ЇN�'�DY�0�fyb���m}+��yUXP:Z���J��@~NX0��&�R��� �σ��k��>�}IGߋ��QG����CjϠ�����<>P����Ϥ)zQ4����6O�R�����qO\��(��I|�������~��Ն�̳Y��\��#���g:P$��P|	�u��%ZnXM�pH���8BH�|�	�"���7�	E���S��cqL��~�K�߬��@�BL�J�7�R�,CD�دj�y�:	�	�G�Oh�J��߫��M�ԯx6��NW�v��R��[ځ�#uጪ���{����X0M%�.��]۳@��i����ߙ��릈�eu������(L)�x1�:����+Qc��`���I�oPd�Y��7[��^�4rɒQ���	�:@�["�B��̴R�ԈAD��Fw�`w1e�	������ꗒ�q�b!��4���4
�`o��^VY�Ei2�w����݋-4�(ټ�(�x]���pǶCB^ԓ�`��ժ:at�K"��N'y���)�b�)_��q2*'L��z�'z��*����X.|����X8sq**Uq�p�H#C/�&�o]��~㵪�l鞪��j�]5P[���Kh[�]G����m'��C���p�f'��ͻ�ʠ���A#��4��&d���z�]r���H	5G�^y���q0�������������3o��U�xׇm�l�|�&�LJ�����؟6�� �UDg ���u�L�j&潽(�X J�$���یj�d#*�VAb�2�Dw'�k����4�i�]���|�T��[*Ҭ�)���_�U��0�����1�i�<�Ū旴��2lOG�ٷ�3	~G8���"z0��&\kb�ݗ�)�4�,Sjd>���M��h�_~ύ��VC�T�1�<�B��A��%����3f��$��94E62�Ź�]�K^VH+ӭ�j	v�A)8��q����]���!Kf�j-���������ȃ>����xkj�y�-zl�x�~�l�\
M��/�����Ѻ��B���je����q��!�o��͛���Ps��=����o����;+QnmM���
5�̘V�,"���;7� �3R^��aG�e�_�*�ʹ��e�[:�sw�@qy��Q��c�M���S�Kw��Tns�Lm���{�X���TЯ�p�?Ni��f�|u�;
�x媴�F%��5)+f�h�ۏ��y���
��u>uc#�=:�RYw��C��֥za�Fa�������\������.m����[�.��=��r~ze��s�S��}��k����1��@��j���1���9�ǈ�SInV<�oI| D:q
�Sc�� @�$�us�q,�Vf�_�ɼ1���p,��+ �w�s�ӕ	�2s\���e�.��<�W�N��*n[|�˝R���Ҥ,�P��v�F  �
�m�SL{\�4*x���^uwzQt�G��c$T�������jV��s�h(�Áp~
���[缍T�����������4�c�÷3fK�ln�z�H*��� �nr�R���ځ�כ@�Co�iv�����Z���jI�31��w��v
A����;�/å|�x����4��2�Ě��2���C)�ӧ��9R?�}{�߶�����~y9E��"�ݸk&�Z��QrIlba*���F���i E9���xSu����N�Um�T���lM�':��,��v�1�5��&|���7��5|�/8h�8��3f%4�wq.���ʰ���J��>���Kԗ݋�����<`�K��z�6��t-����@�{FЀ&bx��;�I�ƕ��z�vGu��� � Y8�$t���� ��i�f�y��]6䪣��[;X��]����7��(��z���>����o
�uG�A-����޺�]J_i��_����p��.��������Ir

(����9�X��&���m}%��u��k5>π^����7�k����rBA�!��.� ��\�5{p������k��["��˶%L嬌�z��c�$�3�>���g�Ӈf���F��O�=I[�2-�0��m��?a]���D9�<b 4��ޜ��L&�Eu��[�u���I\�S�x[.Y�жg�8f��w�1���]#���!�'X����v
�xL�"S7B�5��z�B��H�B���'���y��RJa��5U��x��z~ӴШ-S�3��ܯ�K�VZ'��~����I��%s��nN|Q�cTm�s��#�7�T0%�[P:�B`�E#�*�ʏ�:�W�	�W�����zI��ǌ�0A3��!y�)km��Z'�u���v�'��i�ޅ3�_<^DBՋ�kA�n��)�@o^�W����ʠ_�OU㧰r�4֠��q˒x��?����X/͠���=��ެ�z~���i��.z�Dd6��W��ӝ�$	s��`̀H�وk��	Fhc��Tw��z�_�5*�y������N���fo5?��@�:�/��������2�˛���t;���ɰ!S��Y�q'�
�����*-E�����qM����S�tD� �	����>�]�LՎ֎�(����+�K�e��e(��A?���/O©'$����~]:SR���[�8�y�4,�:ܓ|_e���������#e@�R���Ѹ����BO�쎯o �/w��I���,\W���T�Dƛ�G��i��LK�`<�h��W^�5ؒ��x�6�x����IҘa{!?��@P^w����.����J���Ζ���M�]���5�YׂUث���A�p��� �l*�}Eɰ,��;�-C���hv����=�w�<�8ס\j?Gd����z����N]s�O
����l��h�)>]V�� [�����p��xް����ý ƕ�v��	��DA@��|�j��QQ����s�׍��s�4�̼MZץ�_�
.忶�X���Tؚ�,�#l��μu��o:P�D����'�q!�����M;�'M�����(Z}�"a�A���(`M��y��Q� Z�;)J]d� z�[�^N�Ȇ7�-�y���֏۟�}p�E�k����Mpx���0]m���=��"�����?f��\����6�`H�Un�q�Ka��Fă�C˧�k��L|�<�}-��tV�+5~����>e��ν��5��>}�ݓ!$�fR�ٱnXe{uz�T�px�p�x���z/ӟ���u�R(��J	ds��������7`����� Ն�Z�H/B�Y�6Wh�� ��(��A7�w��c샌��|V��� �ޟ��8�N���Z����Ƿ$�*���M�@�1��{Oa�Y�r�!ms�O΀z��ٔ��g$;'����Tު?��y�_u������ȱ���s�_,c�ĸ��O��&�\.�`��W����Z�Q�^g�Է����Y�ۍ�-;o܉FFF8�m��&�`���MK��a����r�=� sl+Uי�~��O�*�0ί3���F�������{fW�����-�w�H��<U�d���LVIl�!\��ϔ)G]�]Dő?��h�w��i_OQ��E�n�X~2<?�c���q;�d�{���vh�ӥ~��=�%ߴ���Rw�[����V{��" 	N�«w��H`��6�8{�z$ ��J@A/��G�^��j݁)��bҊ^
$��$��TS$�ַҼ��@��Gݱ�C��ց�F&ř��w���8g04����"d��6�N�Y���1+c&Kp�!0�t���M6��/�w����������s��>�}z�,���d�J�^ ���/],��9�D��KQ(T�W���K�N7��t�T:N<K\��;k��S� I �Nu��k;�QSx�:=�ˣZ%*����Jk����r�b��7a/�X=��l.M(^��g�?7�?FX 0�	eW6'kџ:?R�����l]��́�< �2�2���Ϭ�gsJBBց���R��vrR���)xKƴ�u��K��31�<s�:4JS�'~�4@�i���ԥ>́��dL4^U Y��ڍ|�{��w1[��t$��(�^r3�e�D����Ⱥ���sP� �S� �.�+G2۷�ئ ���m���@:�3쁈���tS�>'�o����_T/��m�C2��1|0g����a�~�K�/P4�,��|=$G75� w�FV-gx��2��hTp*.̑�����E,T4����+B8�x��	~4�Jwx��%���#�Q/h�!" ��r�D���@6�PҸ&�H0+:G��4 n�Dm�NQg��?���U�:P+:jF0,xBJIY���.O���-���M���p��Z��1!ӿ|J�mIsg�J�ʲ���侪+���e� ʘI$zS4�p�+g�C�S�y��
0b��i+�k�F����a�K�ʁ ��1��#�Q��V+�b��W ��}���;\�gɲ�R�����^�k�pB�y�����ቇ�d�M�X�U��q���k%I�&βS.���(O8�<^ŠK���j����1�RDm8�$\O�.�*`�؅��W�%����t
 }4���4�X�� �������H��������Շ�;V��|���:+iw��@�5u�E�+R�"�N���y�?�>�o ��]�3�ń��$���u9Xg� eS�.�0i��	ϝHy s�5�U[�Xց���� �YnXqv���w	n�{Vp�t=b���������˫����M���I e�B+e�},�	��Bs<�(���1��/E�L!d=�%;?��Dα�Tחp�-�!����C7���+0�[cr0�%�J	WK�EU1�n�>��&om��"5�hQ��g��(\�����.��
�w�5$�+غXP�3�s�n�4�V�!g�M�~D�����܅���E�}�y��[�/s)�V�4��u̴B�I���&٭�e���c�S�k
y�u(`�z�2�+�VE�1�OͷP�����6pf����*�v �@ƸΫ��74��ߍ"�&����/��`�����A��eP�*8N�����s��Iq�X�$z���M3���}Y��$��$�x��
썡�|�|���R'�� �e[����Z����z�,�m�q*�n�ݚ_� �?:3�Ӊ������C0Z[��V"��o���F��	,L��Xs�0�,��h�*y��RR���]9IH߽
RI����)�}�5?��9ݪ�$\�L���2r��� �{���VՒ���*���궋��m3ކ��G�H@n�dY�0%��)&��6�Q�n��Hѻ����k~ۅiT���|:L�P&��U�o�4ێXHU�^���TS���zÚ�W���继TOX��Z���Y��,:m��yU_J��	����r���z�?�x]��ZL��T߫@%�N�O~E�r�>�V����^�!��U1�h�À����7�ƦO��Pʊa��N�%;���}]AG=��Zk�tt�?�u$�(�ƱYZ�W&Eo����^O�.{�U�W8�5�ohͲƲ`�k�gn��)�QDA�.�ʌ����?��ye�\ 8	H	�֋�Vl,WH��6���;��)1@)
�����.@*@���4C[HSj^�t�K�,gS(��h� �t���W��Lz�:�{� -s�Y:����ө�tD.Ѯ���ۄn}�2��)Ų~K��#�D����<ҢeZ�%��cD���g�KD���5��^��XNq����������Զ�s�����1iv#�Bd|Q�4z��[�p������|�w�=}��6�$��c� �`�#wь�M�M���I�&�%��>d����'1s�v�*��}w$#����L!\�y���a�fHJ��e��8� �4 ]Cؑ!��x��c� |�i\!�-��yq�V��8��c�5H� xJW���W����ܖR�@�H.����p�,�u�)� ����K���1Ў᪻���\��]QV�ROˁ���s	�&�)4��k�����ĸ��D�rh�\ӟR���ћ��y]HvJ 08��|I��jnÙY�`��!^s�`�ߑ]�����l�"��S�d��`�B�`�KXq�����@B7��riYr�?f��)ٌ3�Ԯ���XC'�k rV�K2�0S���o �ڒ����ma�k���F���&�EM��x��u��Z"��*��2�@z��������F�<'�Ȋ.}ߒ��U�<����`��P�����V��8�3��؜���#N;�>[t^M��yv�\Č�u�<]��4��o��>�6�����yd���;f�y�7E�c�)7u�䌰j��͌7���Q�z�-6t�?u���B鶴UŬY�j��ec "�^�Q�O�Tد&�e�����b�Z=�!�i~��-�k��`�	��Gӽ���!����bL��3z���������`�Q,�V�@ �J���������e\ø~>�Q b�D]�	�l`8�&/�����FqA�٦C�0�Έ]Z��:G�,�`�ȳ4Q\B�mΎ�]{ Y|'�M�R�]}��ЗK���Nu��x��AB�W��XH���D��<�Y1/��*N�d �UH�8|$�z�!t�|��v���XG��q�үRQ�&�R`��$1�t'��]�1��UMaF|b��1�(~
���5z�ӹȷ�g�Κf���m�\P�c���>�gGx��YU'��5B�����;q�^R}{������2�f+N�`c|~�W�j��?�˽�3�[p�H9y'G�k»!����ـT�鼕v�Oj��ߕ�9�"՟ m���E<ie�ȢV9۝#+�C7$R�T����)���YYL�d%nWbo�s���v��b��.�;-�J�(��	^/6	���{K{�$�׬p<I�����c��&S���s�:�m�@쐅�����i�t�wn��]Z�^����{h��r�Oh��)s�S�x��a)��<�{�Gހ2��pD�fIu��Н�Fw�ͳ�j�r?$0#I6�6��~D�F
�؞��꺠?����i�zw�8"�׮fO��W���ڤ���M��V���Z�W���bҩ溧k�~��܇�;��@�h�O8���ϑ���!�f@\~ٝ���EH��u�>�v���Z�J��R��E����Y	���SW�Ƹ���T��-�#�������C>6�}�?�{)��t��Ww2�Й�x��4�!�g��3��sw8�/.�K�k�D�=UAYˤ%���>Qz{���S<l�M��ga�u4�d�]~w͡m�E|P��3�?�E�����v.�?߷7Y-��6\R'��d^nmɋܚM��{�ϣ�n=�H1g.�b�uޡ��,�ӥ�P�m��QK2PJm�Uu;0"k�Kw�Ӣ�Ɠ���n�<dC��ml'r�~Z�Lݰ�C�ko�V� �`�c��T�v�#�D��p�8�=��yS�V���t$�틗S�u ���1�̼��o��D�;4r�IXQ�-�)�n|X�m�{����X���m�Q⓪�fc� �y�i�Jߡ:�^����H(&"���:P��AU�t��B���0�~�6�WPp�K�.ǳ��}�=�TA����hg���3�B��U�mN�P(q��hhŚ��A�(��QW�s�.hY'���9,lg�J�CP�'N����N�1��⦗յeX�S�� #W|��X�];�����/�k5+����
$PnJȢ*C�n:��]D�؛����5N&������gH��N�r��4�@HUom�19q�dTU���;-�W&5��~/Y)	҉�-_��!���DRtZ��W�b��d3�9��ڏ�\�~�� @�H�}��v6�q}z�L�a���6�2H���-��]R�r`��ʅ��*3��N�1t7Cfgj�p������K����ծ�h-$�<�{�+-ڻ�'�/�Px��/��7��0_?�u�-�\!����9���d E׈��'SP(y�B�� �[��!��'/꿬�M��Z �H��u�$�E��sI[�"�,HG���uH�D~�Jmu7���U�6�����*��f+N�M���i��w@�I��3�DÆ1g��ɑM�C��8�����C =������.�0�m*�/d�`�����Ԑ���Ҕ�y2�R��I��C��(&gZ�+���E0��y�7�x(��:�j�3P��T|��*9�N�)���Q�gH^�|ϱ�1��ffX�B�����G�77o�E_��s��<R�i��>Yp��v)���c�8Jm�ԓS�׎�t$�h��SqU<��xiM�(n��.޼1�~ T��I�d,Q�Q�B���oCsK���<Iǉd1�p�#v/Ӕ*�*7���9�0����LV� �}a3�R���&W	x4)�}7�h-�*���Kʮ�v{��zܖ�9��X?��o�t�����ic��W�Fuҕ���d|��d��b�{��^m�����u?ÈJ<� ��\?P��H��մeL29夢�S)�-��۟l�)�c�k�R0oQO����9���?e���;�_ޔ�c�Vy�,�~� t�vo;>ݷ+_�������K�/�V�#ޮ.��~%G��N���6��O�N%`���7�DD�b:!Ž��p��tӻ3ٻJ�y��s^�(���h�p��Y��A-	;��N�}I��!�Z^�M��u(~]�b���?��ܤ2��_|�l���thjU��ſ>_�-2-R��e�a7&��ũ �o�%9_����Dn/��-_n�i�K�י͛h�m�G���<P��7�hlR)��#��.�^��Y=�x��q���(����R_ב�xN���9�im�"۝��Io��Ĝ�q��&r��ʍc���} ������!�������\|�a$�2H�/2b�Y��]��	_�!L���*�1�m�[�(]"��1�=RM����樂���՚5���{�j��Y�d`)��@l����{O�:�:�����=D#�ޡ5X Xq�����}I`���S��m��Nz૤Fػ-�/�_�j%��/26;��S���4���~��m�7m�ma3?�-]"�GM=u��Ⅰ\bܷa��Ys����@[���?��N 0D��p3�E��ك�5�mf>g2�tM�~�TQ����9M�HE�i'<��<7����/���j5@s&���t
� j
�&���Oh
z�������γpЦnl���n`�m��i ��%)�	;I/����-���oz��\��3O���;��E���S��g9,/e�Y
�O9��S`8P��xm|�.���xɺ�G�nsY;����w_kMIi���)�W3L���tB�cpF��au�n+� �bU1��-��C�hM˴��ꀛ�%��$"�g�a-�`��K�Al$-�a������q����+|:x�������Ѧ��TN��r���y��in����{����gXG����)�}�R�\�<�W_\�_��xb��f>eސ�jc����X�v$ 3d)v�����uU��zas��bAWͳ�K\r���I��v���W�Ӳ��0Bc�o��7��2.����<�\����P����{򺯕o[�AԕN0XO6	���o����ZYX�j�E%���~oF>��ص��fֵ�n�F��Au}�~��*i���r���	(�\sn0�͍�Dl�*������EV}Xo�`<�{7�az� ��"�`��Az�#�<��gA��#4�^g�	2��]���
�����v�<(f�Hj��.$Q$v�4D���j�Ta��3�e�jp�8��W��Uw\t<$��&T�����d5]XT��f|�궍2k�o�Ϯ��69,T����U�<�����\ۤ�R*��B�x�M�y[xT*���{���BZ,&�R���;G���\F.�0� ^{�5���U�y�X��I&!���|�֝�Fq��ѯS?�~\�
���r�"�0��8i���&�{T:�f�'�Dv(�)���X��;:Sr�+�'爸I��Bm��~��7�r3B`�E�������j�&�&r?�E�>8��o�sG�������4Z�Fg�@ע����p�/�01dcS�$���_v��x���܆��ry��I+�A�q8���Z����f��V,�&�_:���g�A�Ϝ�iT���e'I��UB7����n�?�rM�-���G�OL���ct	dDW����@@S��ž?��U�oD4�4L{�Ypg²>��4��ý��}��:��Ⱥ`�s����1���&�����<hny��'�s8�]BR�h_}ɴ8݉e aJ���]-���y{a�M�Yt�~}�R�0�sE�������Br8b�D[��A}���zj���B� c�k�lB�ԭ��S,W]Z��?�+����� �|�9dt��IA�
��׺2 ����ohf�[ ʃJ��b��#õI��md$��REyx��	1�v]�n��x��m�a_K���e�-	�:�W7GV�Z$	�o[ˀL�a�把�,.4>\Q�ֿ ���5,��/�^��D��ͧ4�fClb���UrD����R�,�I�әtYy�
ӅG��� S�Qק(v@v��s���_����7k��Y�'���
r��B����x�	� &ƹx���/u��v������_��`ߓ*���߂���#������b�H]� �i]t��r0������1pA��Oc;6O2�T�-��De��E��(���mY�ړ��;�V�5c7ɀ�~_ ��j���G��ŶKsQ����\�-���U�pc ��]�La�^MW��_���w��gD �0;��̺�B��u�dm-ßl�8�kK�kvl������K̶�c2mخWɱ���`Bo��s�{W�rV֭~~��wg�:���,�$U^��&a}�L-n�R�M��:��iऻ=�( ۃx��[���	�4�u�-"���Sh�������7�v��F�A���_"��a�"�=����5���U��nL��`�*U�K��4��Y���h���^r�v��eʍ�!6^0~9���F��{ճᘻO<�����=��n�ǡ�Q
֨����H"ZN!y���d�#���dP]ٛ��kT�	_@>A���)�&��`?�1>|lh�CQ��)�y�E"\��ÿ�(��Z��#w�� q�n�I�a��I��d��pK5�"�ÚLE��c�E��P�=�Ϩ��iJ�0{�z��b�[H��Τ��d�u��_�{i|�����a�uvUe�.X�����>+V��B�t����4�40
�m�ym( S�,�=� �3��7|d��o�+uxW3a9��9�����f1�n�"���$��(6Κ�.�U|N����j��r[�����$M�X����H���J@��Ʊ�T6�O�R���L���\�N}톘�M� 2�N�S��'�ug��@#� v�Nm7>C�ٞ�)a�&��=�*Ӥ3�G�,_-N0�F*9��J�@��▓uA�K�G�@���K݉�:p�L�[�M�}ɬH�^5x�G*�v�H�.�ల�h��HKK����B�"�;DL^�l�(^�"���cMBr�� ��J�vs�Ǝ�#�`&@�?�?EN�u�H����L�!��nnٶV���xO��d@W1����lfA�q
gǻ�U��/	�t$X�����L!if*�^�@.���,/p�L��tq"���l�l�K��8�Z�y��qB�&|�H"���T��S�a
W_��G3�K��-YTVc��Q��C�>�o�c��v쀄�N��R�H�Q���8��9,FU���e��{�^�`��W6�粼�Wx�=R�N:���/��5+��T��1���{�_Th���J�YOa	:�B������%��/K���f-�eÃl�F�������3W�uWZ{�qϞq�5�Ua7I��YA���~�?й�d�!�Q���nP�<�و��&a�^�ĵ"���y���Ҵ�dh
ɥh3}Rh��gߍ��>��-75+���f]����FI�k�pPf��b��1��E��+�&#bno}r�!����N�0;�;AA[�Q��s��������]��vQU��S���y0�W���	���BgO$d�Z�-)C`�1�С�qS���_C��k�� ͨ�	�	纑�c����yԊ"#� ��}��cCm�,��(ZfvVw�/��V�m����Y�i�=ы�Ȉ�_k��ٮ&��`��;���)k	�`�|g�Cٌ�����pU-ew®���B�b�c�n�@�3�9��z��x�U����O%���K=U�>;,J-/�j�g��|T]���0�EmC�W"�_^��{�OІR5�!6P�X�u�0�n��9��6��Q�iUF!@��D}����Χ�t:�/U��4�y�<I�"��8I�Z���� �`z��WՍ�#P� �<���c�Q�з
`�5<�|�)f�J��C�>a��ڶa��4�u�h���XŊb W�vY�OK�����[����Y9�"�BZ�R߭7ʫQ��W� 5y^�پ��Q%^",6�:��'�����ԯYBY�6a\a���1h��i=��q	w��@�-��A7�%�=��yl$��gd]Q�EfA���	�ĚY�f��<�ݼ����Z��R�@*�ٿ�C�z�x]�*���p��P@t�HsCZ�i��E�o�����2 ��о���(&�C�w�cȨ�.��@�n��TX� ~�qx�r	�_�,IE�0/�/#=W�W���<��a9�qi�����G�7��c���=�&�?�v�jx�N���5����
a±t�w��9��SS�� >�������H,�2X����;����ۣ��N~&�H��RI���H�lv��p��	���n׌9��f�����ǣ/�-�Ɔ��w��#Ì�S��S��/��pe{;F�⨁,jc`����6;X[9V�[��4��r���N?�G���?�L.�]�����J�^P�a�/�̐_�nK�%��PڶS�֡a�`��{q�B���η�\m9�P9by����:�'��9�<|t.ݱ�nyH���֎��h��A�����PbjE��#���h>�Hn��S1�تYԌ�N�^��2h�B�Q�t�doM[(��ԩ�$�����Z��;��O@���{��̮!����C�m����
�=����3��k��%�ǂ�WP����Buۏw�L^Bʂs=�	JHvw7�^�HE+��0��\ D��yv�->�q�Jw2��Q�_~�[�v�wb�oV[�!�9Rʢ�7 ԫ��X����n�2�*7��K���.�J7��"F��V��s��\�Ld�טgJ�[�J�;_�7���¦� q5�̭F�dW'�=�8��)���#�{<n��i;��?a�~.�؇��n4��gо���MN��545��v�ҏ�R�-(YU�a��p�1��Q��N��%��7+���A���=��[H���.B�OIq���L0�r��S�/�[b���Mסgg�P�eo���YN�@yO�芞k�1��^/�O*|��P�M�-��@9Tu#��aR媕-�h�}:sZ|u���`�F�K��{��TyS�z�}�M�;uZ��"�W�+J:lɕt�:��)N�@io
�cV��!�������HI�0�墆,w�+�f���b�o�u&ܗCi�e
S��Q<T�Y:���Y6
��Л�9��S.�M��v^*';2y����@�=n�{>�j�æ�_;���7+����@;ᛌ=��k�� Lu�$���%c(F}��F��Wע����M�@4��ٺ<���-B.�ټ��5�e�pYO#�|R6��E����U�)�K����F�t��O������Z�9.��=Yէ�;G�x�,v�h����xC��)��D3��/�������r|�v��#���e�I�)�])X5�q���I�^S܈�ٗ����?旀~��7��Az�����86׭R8s� �P�6������UG��0��䓠S�k6]���J��E�\Z7���b�-�Ɵ��5�8�-��1���e@�Ŕp�Z��.�[�g{�t���&����N���b���Otq�m���i�����(�BI�C�t�lp+�e/fz�����V�/������Z=u���I�y����d��A�s��#��_�F`��I�g��|�y�c��.����;N�4m-V����2��(�����mJ���}�A�CS�����S�T��w�
zc��a�n���/���Hk�k|(&nݪ�v��+=h�d_����&��l8��_�t`&�������N1���)5x������7�̱�G	v��3�B�8�º��d8�	���D~��8�^t����F}E´N� sHBF��˾t��AI��>�D%���`��`�������.����v�{�I��l�����V5���/d�W��_����0\���~a���h�����m�I��U�)F��A��V�Ժ����j
Ⱥ:qQ�Y�F�7e�z)������K̇yYϺ�m�vA��s2]�. �oZ1m:��x�����>9�uG4�H+/%�N����7s�O�7
u�,��n����>"��{FULS{�ԅ9��oJD/�"A��f�%�i�6��^����\F^� :<��F��T���ʾ?���<���H���G@~/�q�^'�_�mWH,�Od���킝�R��z��c�c��r7W��T.���/XL����B�	��U	��1(��*8�`��h@�. ���'�5@Y̜L��i�;Є���}]X�5��.��¼7#�d�T2!�]��w2��9�:��ӗ�w��fJ���a�
��;"G-�&�> �_�OD�N2���ϵ�hNT\�#�D?����1�2Ƴ.�_� �&�N�B��n�wޯ��(�	S�.e���Wu��N��h3e؇�M�	�X�ŤM��%ʵ������N����}(P::8
�Ǟ��v���i�ۓWP�3��Xj0T�	�6+܍3y�adF��`pwv��[�Z� s�q��;o8Ӆ��_+�W+�|5�����A�XxTӅ���\�L&����W����y��+����M��3�nH�	Nc�<>��]��>��	V�m?p�M�J���v�6��g?�$�i�`.Q����y6�~���KHAS��(rW��@- [���r�"��1p~�FDa��0�Z.k�U�����J����]Y�y�j�ȱ����R��F����P�s,�Kh��=������[)5(r9����lѣ����-\��dyw^}e���?�ud�7L �;��=@W;e��@
�<m3c���t{��"e����ӒR�EU�I=�q�3�P���O��޿q��kk�z"���:���v��DLJ_tJ��sRs�b�v�/b�|�&�ޱ��zP(�<������D�)�4]�S�Hb�+)t��2�����|f��a	ț�v\�iSm2+��{6<�O4f5��,h1D�o�q�&A&���Ҫ���sB�=�;%zT��xS�)ë�����e$�T�zkz���NV��@^[�O��ة��Oh����I��W�훐��p�vk����kX���AV�іO���2I�*�3���u:$�d:&-�PE�~Xa���(!����1�}�G��})�:m:�9�Ŏ{�yM���R�����Vl^@go8����6�AZ�1�y��E�p�P�OH��:8�{�)�ޡrPD�{(~}�G�?�k�w_<	�fr/ꪞ�I��H~�(��sh��~���"��#<p% t|���o2n���{e7��KΩ�0׊�7OF"�E��ts�l�g>���ϵўT�7�E�+w���O��b�)L�a�k[W�d�wk�s�(Kp7Dp�4��k�ʔ�;T�I��^0����mF�Vذ��Gmn:���������@�N�1�vS���@V�]���ކ2���ؐ\�,���:�r3���ѓ[	��]P��#����~��d����/�����c2�-2j�B����n�cZ񀄄�A�¤��.�C���u?E;7�AM�M�;���+}���򫴝='�Z��Vf��"�$�O�W�-l��SR�=�\U�q���U�(㍻_�!ܭh[�%��sU��y���F�OiN�A�������/B8$1Ф��_��FH ��}D2�W<��l2�;X� �y��/$��&�z,���CՓG�%f���Y��(���	h�"5�"����$F
��{VԜ��f���~s�3�OC�&~���7~���p�������6:��A3�l9�Z�3�Ո6�iso�G|R���C@XHGc���J�Q�-��e��� ������f~�>7��N!�O�Iu������?�dT�u��z�\�#10+�̎Ǣ,?,+�}��)VB	$���YE���梲�����;\ F�ԫbc��sn^ga�Vܝ�����|u/ӝ�q�s���+#�]'8��ǅ$P!8�	㈑y~&��sȖd�*�yY�ԝ��jV�����o��"bM�"�[*ߧ��ڮ�B��~�r�������E�MX:�l�s�T��}���x$�ȭ�7�8+��x�K�pC�r����H��v+�n��t�B�k�ΥN�4�u�C�	 _��wpS<n��X4|Q�_�#t53�Cw�%�Y/�<-.��H�B;w�'���Q.���hO�v�eE|�����`�%�,�N�� ��,�+�G$
A�@����ŗ��{z��RAB�.N�?8s�q��ri4\����_�����1�߲��������uTeW[>�b�V�j^�&�G�ʖា"f��R�4&����$sZ8�w�Ho�_�NM.�^bR㞘P�MjO���	�힝-^�����ؓۧh�,fY)�[��L3� A,v����x����d�>b��~*��	�v��>F�/����qL���T�k_��j����*se����3�g�L�S0����sUd]�}#����ⅺ���-�#���cG�nn�A�z�P���z�� "�$߾��\�L.���a.7���p�NM�x]���r�[y?�]�K ޡ�
m)�k�7���ê��d1�вQ���j�&X��m�f����;Y���nU�^�,0�扼t�e����(�+��g�5;q	*��<i�6۾��]�ݍZ�M�z.��E:���n��2�W�x�k�`�Aj�[J	�:"�tM���՝������2���`���E�(S��OPfL�A�JR~�ӥD`�[~��s��|���$��P�lTc���]K�«<�dǖ�+I�t����n9Ú��7�9���HG2|�=o�c�Hi�t�;�HM�Ʈ*q�*��ƙ�����H
�ɵ2�؀�\�d�S2].<>6ԓN�6%#+-��ξ��#KI��,S�����?�����6��j^��{Q_����B~���w>ϼ�x��ر*f�Խ?�Y	�"����
���pAu!������X���U'�I	���Csi?�8��ۑ�+Oqo�EQ�������f�8�_��,�5�9d����鸮�Q?��;�4��0e2}j �_�0��p��[+���5Ѯ�w��s[O%R�_��@2�bC���")�!��U�����j�C���a��Zw�lܻ��I��*���s
��Bz'�
Wk���GF=޶�qWzs��Ի~��9��?�Y��C��gl����T�~fJa��k�d?��uj��'�.[<�9S���Fn����D%�<��n@և���/�z�����Y4�}�g�>FwC)���GC���B�ڰ�<��sޘaNs�ƶj��,t�OG�6�b:�z�X��B��Ve(B��B�kW�c�L���YB~r���wKk��.�m����r���piV�3��K���q�t�!��t�D"���L�˩��β���KӢ4l���CG����L�:vU׀į9'X���� 7v�Jf�(��0�6�7��zޚ�/̻���5�9wO<|�<����(��P���i���lN�yܣ+�ҏ��L51}�o5��,�:��V�X�ha���B�&�ϴ�m�1�Y�`N��N�`
�>��
��X�خ[׿S���+�*f��� /E�6���k�a�Tȗ ܂��G��ۤ�!��S��U�����3��"j`WIs�4��9Q� �;5�U��r#��R�g�8)l��+�)��] !
��{&�^�8ڌ���
Ћ��:h?��2��n��t|����m�,�a̭-��j~�,�?�C�8r��(n����)�.�ja�j��a��S�y�z�7<�W�g���*4�v2���Z�l��Ǫ���W�5#�i�C�@ƚC��i��O��;�[̼a^�����0H���h�{JL��%Ӌ�*�p!��N
ˌ 7��
p'E��;���w�����9��^��IL��dKwٱE�V+�[�-�0O*��������ҙ�Lj{���'p:������U��������ʊХ'�$~�j_�cp@%C��L[T��V�8���Zd�ܒs�p?b}��q{�Ad������P�y��?�pt2+c��|�d�Pݹ�'`y��M��J�T~�_{ژ�غ2�\f�6ZK3b3_	TO9�۞7�@%�?�To�T�Y�œ��w�w{�LU>�Z�.��:� gmn\%p8�}Տ������A`%�w��dɬ(]�T��!�6YRn�)9Xn�ਖ਼kK����'�N;%��oK؃�!oi���Q:L5HS-䲔J:������y��6p*b�6i�+����sc��9-e0��7�������I�2�^3�Ve�����:��^3�j-��<��[�ꈏ|<8k�]A�� F�+xG�*KI3����^�=�Pzɠ$����l�&mkM5=�J"�߼^V�ɸ@�9�9���aC��®?��)\#���]'@7���9��|U����Z?S	
%��
�{�$�W`�åo�P�L$-�rC�8x��HAm�7�U��j�ExAI���u�Y�B�F��pX���b�V�>0��o�P���wo*O�;d�_4�T#�/f)�;d��:��*CksF��LXT�Zh�M �<U����V��s'����9�W�,���{B��[*DA��OJ(�+��s��6Nf<��n�}<^Ղǂn�ԭ��-�*>&t0�%v�I�mÁ�;��$vL�7�1ӌ�Ɇ��d�X
7j�W��}��uõ]9��i�s�[�� Y��M�4���������F~,�<��V�.���A�r��p�I��V\n)
&k�����l2z��i'X3�E'�d�VU!�=@K�펃�E��P ׀cȭ�����CdВ���*\�h PP�l!��4��S4�k�;��4 �I����#U�O�.]�O��M�.y& � 7mT'��w� 펝�7EV�� ��VeuBӬ�t6���l�ʺ�tGQ�c"�������n;pw��ˈ@VT`Xn��2ϠX�_^ڋ:߲�!m4�zq}�{�vB�_[@ rXF��9*=�w*�mf��v1*���9�>�O�
SkXӗ:��$tE��(��R
��X�!���;^y!9���ȯ��L�x�ƳI��e��*CD/s�Rw��mE���c���g���6�ȯ	!��ek#��f9�}9ǉ�rg�>�!
<�F���A�>l�>��(;j�qE�� �߈aa"˲�˭:�h���a>��	�6w3�����ٜ��:�K;����F+�9e�.�P��I�%��ذ��l�y�![x-����-��w���-�߄H��qږ*V�k>��
^�UF4Z�dvfη�
��hؤ6�7�TΎ�@x5�\�ӏb$Zl�yߣ	�����r~$'�|t��$ ��z�?��ی��DR��u\}SG7��m�*��GΠ[:��U�e��e���������_O-l�SWjJuE��Չ?ib�7�e;!%Rv�[BŐ�,�o��z1{+[�;g��فwԠ.�+j�ߪ�1e�`p�ъf(�"���g��M�0/ՌO�d��S��" �~�&~�Q�<�럲C�U�JB�Ց+�b�h
>��U�J4Wߩ�C鯒��9���F1W(%W�$nR�&�c��������Y_-�F
0~�cy�k��qZÂ���� :4��\mZ�F+O��p��`(�i�1]ze�RQ�8G,��3�	�s ���q��$tƵ�9��s
�G5��O�$_�F�7��"��B~�pk�{��_�����r�T |:��9pJӆ��
c)����
�k��7w��&��yfb6�3�c����19�,����';h�\�c�Y s'�C���h��̆D��?�j$�^� ���Q��Y�d���<q0�74P4�͖T�	���V�����݃9���YD�ihᶤ��H._�Cɱ����g���=B�{��'p���rj�����3�kV9(Y@,�Sm[ߙ��7)Pq;�j�M/Z�wq����ћ�YR2 [^,p�6 `Š�'�q�R�E�S��y8\�5�<v�bQ�1�O[��N�]�ŶS��m0�<�3،,vS��+l$	r����Ѩ�� yK�=1��
�l�lU4�r��q���!o�%_���ή��z Qɻ*���O%��Y��r��+\%ԝ�w�T��r����add���B@���xÊ��we����2��h9%�b�� ���n�6�lv���4�����>�O���('L���I����Y7��'���=��(��\�3�s��e� ���>۟���O����+a�(}��i����� �'=����Gd���깅kz�s28��i:�m��"����-@V�(TAv����V2aͤd
���%{da�h�[%34Y'�;�����I��x!y���h�׷je�=>4���D�8��/|��a�B2ɻ�?�ڼG�z��Nϡ~H��S��b|��D/]pT�� ��+��A\����Z<kv�xܷ��|wN��(�W��?��j"���{.�w�<�n�\�u�-�k��&?������������A�9RP�j�UEs�������='4+>��oj�n�d�.��~	ݘ�Ec�?����ޑ���b�"(e�ōU���|^c��Jܨ]T�4}20dy���A�Oǐh ��6��@����B��T�~�&}�v�i�h�fj�~=f���7�͡��E�_=b�ws��c�3�����N�a����Z�-Ed�g'Ƚ)��<:��E��-jޘF�~�o�|õ����ř7L=@ <�h��<�CK�0�M{�X�ZYȔ4}\�V����Ќ��𫋜_/ݕ����Q~ƅ{-:|7	T�?�~
$���7=�F�8�U�����e/��l.��z�G�FP#�Xd� }XD"b��jX"��T6�sH�lT2�d��M�F����[��:��e��ݡ�c?/�R״�=8�f��I���6`�@\���%M�����"���~�����IV%�C�z�\��2�b��0�}dF���j8�|,2՛�N��1�=ϩ.��+�6JI�jR[y���Jap@ ��[�oh��C����җA-�v��W#��	� �7�����B4��L$*�_=�!�lc� ՠJ��5^���������D�+�.X.�D��m�wVF��53R;0E�r�)�Y��9��T���u����������Y>�>z,��2�m�B]QJ�v�Qp ���7ʡ@�ADR���A�B�L�8�G�͠׽5<J4E=�Ʋ�O�� ��#���Yu���$���Ѧ���'��ݙh��Ҝɜ�;��_�J%��{E}�jr����:����Y1[?�Q��:xҰ��]�>Xu��_R{m�%-K��VE��h�K|r"m{�-��2�����'��[�&e�D%���7�1�g�!HZ������[�y��ӹW*�^���[Q����-3uJi{����������'^F1�1	��|���Ю��1\B]6��8(�.��e�$�*�AY�uVil8��?HT/�T8b�8�;�dɌ$�?!`��J��o�t�n�梺�|�T�0"�g�f05v!�b�T�[��U�2��2]�뇭���iyk�N�T���Z��?�_�(0�L�XoV)��B���{(�c3�Y�y��]�=��M�G�D�^)��Y�3���,��MY	��y��G�:~�q�zD�.3Y�+��󤺊9)�\ f{��J�ש }�?-��[�qj���;�G0REiEܥ֫썴�.��QE+�f�6ҥ���` ���YXֆ���&h�)5�%π��6K<�{
~���@E�]�Չ^z�,�1'gV2���#J=����O��?"�4����)K|07)"��e�O�2 1;6Q���ng%pː�b��m��c^j�[1����k��_N�3�؁fX�l��r��X4ʐ3�<��N��D2��Wo�Io����I6C���kwE'�}��X?��0����qNģ�DQ&�9b��n�1��%�[���7�X��LS&���	�"�Rڝ�o�r��7�3:���<�8|[=U��_�E]��w���w����=����f��%�?���<��\�ڱ-k�e��!|����(I7�>j˕$����K�+���PUġ��O�l�]_��U{X���߇-ʞ5o��7�Q1Į����5��<U���k�N1�ĩN|�+�k�?��&�)C�j~<�Ea*�UE+���`�����u�Hd{o�tma�Q.�/;���٣| vIe<!=ќ俑�xX����>9�0�������tm��A+I�u�t�)XW��V�l�e\�Q�fh+��:�Q/��I ;��'��bA��q{�W]F�_�{�x�SchW	�\qI��ЕS[5R��s��K�!�m+^��!�w)�YɕB��{���${����:�ִ��E9�"�e��{n�#^@��a�[�.�ZК2�Vů&���m�sc�`�v�4���0�2Ֆt~�y������2��	3��H������cgF5��NC�Exu�Fۡb~�n��R�?���x$q�ō�j1݇a7r
\�3 �܃6��y�bO쟒�.�e��!�

v�E+ٗ���5�����:�m�6�&A��=��Br2)�`-��H �����' �Ԧ�|��~�X�tf�/��rg$u7x��*���KT�JnM�ai�"ƕ�K��9��)�<Q�;�±n��y6_����h�tx����e��5�˽jtk��C�"�k���|�K;ﱌ�)�k��'��-ou�֠:G"Q���@i�L#i 8^�u}u&�A,���Я���7<61�ޡ+ۓ٩��0�7;p�T !�W2r�}�2�C��q�� �bV8]]P�7�tg%!�Y����ݱs�����X�՝��H�8q��[v5pn�C�HP	wt�{����&��o���B�Y��S�11��+	��CHJ���i��W��+�;7~����,�y��2�`��&������r�1�I�ՄJ���ه�ts�~ƛsH%�l��x�ވ��{	��os���"����=��cy�eN�荘z1��s���Q+��!C����w�s�
�9d�1��@{ZwD���4�p���($T��F�§�w3�w];�Ƭ􉒄2�y��`òj#�`��U�!�F�D���u�J�V�7�_�=� �Ƿ]w����
i��>N�!6hD'P �����Ծ�a�Z�����r���Q�X����En=XA����ɇ��;�K\��-z0� ��>,c���#ʺ	�>#S�QlA�PThj�ty����Q�s[��F,K��r�� fQ�)����h1��yRH���R_e'^�����'��ʓ�ʅA��F�}K�?n�_@*�qS�|��#n�$)�"�h��^E���ȫ����볍:m_WS4h6mD��4�e|`��ĭg�.�`���l������k�X&���1���!�j`�q��C��]jC���2P�,���
M�l!*Ih��\]?fCᛕ��S�IIÕ�)����3Nؗb�� 
��D��Tl����J�+-���������c�T��F4�@Ŏ��W�������u-P4���4��:�~�_�5�s�m�f���8G�Dz�U&���`mb��:���ӎWa��H~��!�����o��x���N�D�mt�L�
T�j��Pvj-Ɓ��k1��ĉb1�gzY������d�O0�\�O�^�~�ʷEn�Z���Y��:Vp�P1���C�Ii$h�]ng���Ga�DXNl�|՝�aK)hԁx�D(Ej������f�d�x����d$.�Ѹ�QhZ�v�@�`��M�Ӝ�/��ۈ�֗B�w��ޏ�ͮٴ��fז�简7u_�� �F���@��þW�����
���`���(�!o��#t!S&���LGx�����$�V1��b����a��?/�~�X�ߜ,Z����׫J|Z�1�$�1�I��K��u�Ab�EN8e�s��ٞq?*3 �����zb��)�C#N�R����eLN�urZY�n<�o�B�����;��WĮ?|�Kx��2hT�O��R�G���4����5S��s0����T8��\x�3%�A�𴯄��Laa�q��+��$�ʸo_��e���)^��A�8|� �I�>>3�����H=bם=G7>m�Յĕ�e�<�G����h�zKH������+��&�M����"*�>�N����޻����@���YT_H)ˍB�@�I{�'��c/���c]�QM��2�A��b���	��f�e*��^�-��~���R\?R��l!��9x'�I3�]Mu0Ut]��»��"�*wp|�p�B%<�Ϋ ɾ9�g�I-��`ZOd�0 ���~��9�J�[C�x��&a1�E�:�A�������>}P���~"k��E�5�5�W��_�}T�7`W��/��R.�H�%}�@fzQ|X�������C6)��*�h8��+)��pI�hGQ��^
���X�O	�!ԯLR�C��5]c��Avg�_�-��r� ����س(-�}�����W$m^q��=Ғ���Œ'�}wk��hx�i}�a4J�O�2m��L�ӣ㢒mGQ��۴{�n��(�m�-���Gﲚ��o��e��W�]֓�q=�ji}q����rj�����������]��:�k�ub�q�%�~���� �l.�t�^�9P�ִ�%�+ӳ-���i�� epܝ���=�fv����j�Fs�#*!-l�I�p�0���	�>����\sJ7�Wmk;�͞'W,��r?��H��*)��-gR��xU�ܦ�Z���V&bX�PI��h�0ܮ�����O;	���G"{<�9�Q(������3Ai̮����c?g�����q����oV�z��z�=�Z�E^}*]Twh&~���O	������y݇��Ĝ�'ap�D�[3��>|<|%��&,����38��\m�PQ��H�k�ͪb�'��̝3���3
	���IZM�j��+ ��Hj�?��w;�l^k\1��g���V�JSj�D�!��@�T��<4�e�6u��wp}r�('��(p�В�:6�����c���j=5[��xq��}`����]����p��y���X��bV:սa��Y*��ɶ��]�5۶�I��E4;9ީ���a30�Se,���꩎�Z��{�1n`O�ԁ�h�I7��sr=��b�G�g�?�f�6�&��0�����(�}���v��]�v$����jͨ��Y`Bؖ��]�vZ�H!X�7�+һ��!��t��t�+�R,�/���CW*��7F -�^@s����=�5n"s�e��CoJ�핪�H�C����˽�T���T��7��:�k�G��$(D�7:��>�8F�~��oj�׺�ꦫؗW;�����|�"Q�	7�ɠA�u�\��1lԺI���'���?�|RI�J�Q�_u�6O_r}�yꘟ]���^�5�_nn&��K�n��u�0�D9��n��@�W�#���ig��_M"�_uQ�@>ŽssY��uNA������g�E����Ę�}����ČCD~��۪����g"���k}}���2�����GB��������켬Ճ�~l��d��8T�<�u�t���ȯ_8���	7=�9i,����<rȻ�#u�ƾ ',7�:_e~�u�=�|��{ĵl�f!ՠ�;9l�MS�B������gzh��GT��ڿ�:2��J��_�.��2Y��ԝ���{F���T:�!`e��&��Yop�}�H�h���gY�qօ�g�4Ak�,�с�r�� A�7���&&s���S�� �#D����l���SM'턈�e����?�|-S��lĜ�SHW���eֿ:!�u��)�9{^���5<PS!U���N�g��ˇ����9�-�*F����y�1>���������P �Yt\9�lj���M=����>obz���@�����t���)]��))��L��)(T��!R�ʥ�BF!��b�L�R��m�@���4W�x!�����N�1uΠ�Y�l�0�24G���W���Dy_Qf	9���Q6��.YCx{��R~�����w�j4]&C� �i��i�B>ϲ�|vfy��U��ڑ�ײު��
���0���ڸ`B�������~�;�d���Vi�$t��z����gVnoQ"]��u.[�-� �Jt뻑��awq�[. H�<�|��S��X����7�歨@����e7�q���"߃sfJ�Eq��(Y�;߭/wn�t��5�'����U!O��T� �t�zv@٨�?u�=���g�EO��W?CQxzN�����i|^i�?�x9®V�Lı��#����B������EXe�9ܠ��q��{ 㿉%�o�q��v�t^������|,����*pkϾ�-e�ʣ�Q<W*N1���|nQ�u�.��)�� �	^'+�	��د�D����tOc�Ȋm�8Hݒ��m0K���Ӵ[�藀}���C�!��絼��i� {�gb���dW�30;K7�xU��)@[�]@�`�6W�g<s�"JlSZ��3���w��z �z�ĐH�q�z$����)1��y璨Oa�:%ʃ�ҿ��`�֝Ȁ�jn�Q�vu#bę��ZJSxx�7SֵY_�z��Zy|֖�����q�}��.��`�֐pvҟT�y������Y� f.v��:pܢ�0�5:;�-�n�L���#��Ϡ��C�@T�����}�5�.k�{ʰ۠/�ٛ��&�b���>��� ����xu��ٓZ�$y
V���x��tApK�87��d#=��bUq����i;��BAz5g���C6�&<T͞��dQf�-ĬF�C���'d��\qԀ
9�2��w��%����`�#�[I��5��3�ev�c7�Lj�G�yD�2�a���P��!B��,��!�:f���O���^����t� ����2.���&�[�E����rT�|�%�H$(�5���u8�h`��D@�� v�r޸��-2
6 [�sƕ�(=� A��=1�t�N4)c�㏬*�\pJ$��Ͳ�Nq��8�3F�#�/�о����P'V4������m��Lto��s�쿟&�����L�w��V?#,�����'1T��Jg ����^���ml���5����WT�e��Cq��E��_\�H+�q`V�.�?�8�~L.��Z�,O!��߄�e
Ґ�f7n�'Vmq���ڄ8�1�R/YaCF��E�#�hxk�ti�ƻ�9�z*�(���q]ft��N�h��	�L��<8��wjA��d�~[�wt�6��$���Ҷ�؛��]4�V�׹��I�f��~E%�M9r$���y*��i%i��Q�摴L:��M��l�S��b�b��q���C�W�yQ�-����_�ƾP�X*_���� ��p����^?QE�y�2��l����eA��?��[k������C�F��=8���*��2�(�lbƁu��y�l�Y,���P�IQS7A��9����f'�ɿf�)��^�	�ȿCh�z]Z�� &}�>�SC��H������-���ȳ���5n���n�����Oe.hd������>p|���5��YX8�xPi 4�OI�M���Lq|*���)� ��!����a�T:�8*G�!PP��ga�ƙ�W��ap:� �6ReH�x���==7�^�>Xw�#�M�X9��Ֆioȓ<wqdL��R�q
�QtO�� ~Q���f���=
�[k���C{N.!+o䞗�]^����!�@�~�#�KUzM�g �5�����9���EU~;�8 �Zm�ݜ۪�偖q2tW�ߛ�Dq려�������!C�HX�#���V|m0|T��\��n�`.}�S�1n^�az�b�lla&b���_%���f��K$�o�w������hnM5>�cl�:M�k��M`�e���r����|O_3�3�@��X�_x�{y&@Hi@h�q�E���h�W���b�)�!�`c��E�L�yq<�Ռ�m�̍qo�=m ���K�KqQ�,�$��a�Gt���|�5<������i5��CeUֈUt�+��S�CH$�ϹH��c+?�r���t�^���6I/,��9��EOsf��`��8�yb��]Ӏ��l`a�na��rUg;2�����Գ��-y ���=3�A�+���	m!g���řؘ�Դ�G�8xk�U��i����pLX�8��t�V�x�!Xف`H�j��ym�W.ZgV W�xEz/��i���;���~�T�Ȝ	f7ހ��1���Mܪ�PQ�U��i1�YɅ������gC��8oql9q���������XT6ٷL�4{E4Ī�y�P�(�e8�����wЂ_���	�#��ay�C �g2Ch��П��������5���isJB���*���&c���Û��c����8��y�"��U���׹}�G�?����X@E����q2�?3[��O�<l�=��5���U�83xo�k*9$C�ةkZSb��U�_��h<��}֕�9��-�����f-40f�~h@�lt:I�7��(!��>_����6Ӧֹ��N��J~͕���R�����{#{N􆃰X�lB��M�V́,Pj�M�pW�o�W����n=#���Y	Y���<"Ug�f����2���zj�/�SM��?��Ӄ	��dr�����8څtgdy#A�bc�5^�"0�$���/g��u���
�� Rh��_p�2O�4��+�D���:����M�?��.yT��4qEt!?�m�w�&.���2�=,%a�9�Fݨ�s[L��T�e���镘#5�b���:*�;C�x�z0�mЋ��NQQ3�&���w�b�`H�P#�����S%�a"�.~˰P��;�)�ةQ�D�EP�S]�;Q����-$UbN�I��X�U�W$S�6�����/�UJ+̝3Z.���Q~�i���w��O��茄�Zg����F����ks�bj�&����4D� �kuqx`���G����<D�s�z	��������V!t�M�F鐲�`~g�j�W��K���e�����d��[��zf�!<.p��?�+�I'�]7���f�X���1<�x)�>�O�q�����WU�|=<Kw-V����_h�Ci���̖@u3�߿:L�1�k�5�� �JW�pҼR~)�>��-p�P	F��[U�e�	��:2�cK���hnS~yMҖ�N�-"e��;.\p֋L�~�_��vl�j���Y����p��ʇ��+�*��ڍT�gB��_� _�A�C�U�Q :�����Օ��5��I���~����'�����RB�Γ�(c��ٗ�o^�E��(d�F�j�sY��cE�M$'��C��SjaƘ��}hvkkK��i����X��!p��4�����!� �f϶ìH�����7��[w���xE��"��p�e�<N;��� Y~�$p���d2A���ߡt�mὑ�_�e��-������6���S����P�m,���[�R�e�rV	�a��Vӂ�Tk��طpn��OUF"\;c�	J���M�����`}n�B����wK�:|!���,f�����28g	�����Ӧ/{����!�=�F!i!ڧ�~�i���g�D�h�ɽ���D�c/��h'����jFda��U#q�2 ;�4y�9������i��X���H��/�Ô�?]>l�Zپ%_p�ԝ�pK����Ő�z�����+�f6�t:s��7[�rN~~����xg8�nN��r��Zm��\��$J�Z�=S-�Uf�&�r��=L)�\��Z>���%��h/i�2�L�P��!�c��)Yd�i��8�
��<>öDRgU4Iy�[�x!X(���F�:�Z��7�4 |z1a�jA����U��5���ǝG-Ԙ߄
 &T1 ,>�d����_�<����e���SF��6"h��Z�ĭy����!�a��PǾ�m���L�t�ȍ�} �-d�j�������ʰ�%��`��'8���C\��/^6x�
�l�����}5���Z�ˮ�ǐ���y`�O����l��*�ǈ؜}9u�~ay]�Pɨ0�]�y�{OɈ���+���JȘ�r&�5o����q�q71�2��k�Dm)U��TQ,�5�X��La�F�f��\�-�Gb�!ڊ,�����`Ǩ)a�<��(p�;���76�"�
Vx��g] =ޞ���c�5�r�r�̬v�~CZf~~�>�l�˴ntԡ��R=$Ч���Ѝ2	1F�C?��Zg���d�el}+�n)�)PȄ�ׯ�!�Γ+)����:_���Z�gX#�Ts݌����y�js�2�S]��.�ru�M�C�>����+�_/� @HA}������Ú��3~S)��Z�yَ�O�|�Q�A�x�����<��^��9iM�ӜLq ��]]�̡n-�I�W�9B/=Z6�<0���W�H��s2��A��bu�K����g��໬���Be��%X9(��k5щ��-��������xD'�r׉8~j���$"�����@��j��+>�k�!N��\���Q���g�@�{�lOJ$w������/?�N������=H��o	5Tn4,�(/��r��8_��z�% z3��on)��"āP0�X[�c�Z�CA%��	P@���;���R���;U@Fc/ݑD�бW���sB��8�q7�J�rn^�Û#[���7]b8��Y����g*7c&��G)�8�Y����n'�p�\�0U��*��3�̸J cK <];��p�ըDf���)ƻ���'Q�?<_�v�Ȓۣ���{��8>�*Y�a��rSI�ӌ�G���5��~��1��%�7ހ������󡈪���3�:��l��x�y�H��k����Z3�#�t-��A�c�Kp�[�WW�c�.	ܹdC���{��W�j�wL����K��N�j���:�W���R�V��x����_�T�E��h�(
�_�za'KI���fR�&�O�ŗ���ϧ���2�6ϲ�[�Y��S����*E��%g��P_F�뺰����^gV�S��h�vU��Q�n)�W�X���gFȸ�K���G4�_{m�&�v�Rʹ:E���w��xf��"y�m����Nɑ���ɧ��z~�A�\S?3�x6j=�l��_<{/����N����ʺ/)�Z48f��M���
��8����4+K�������¹?y�mTg����7� ������y}��$�J�Н�D��k$<I�[��?8�ؒ�ɻД��E���#��H��'o�2����L���?��.r�@O��|ޚ�K�KU���5�],L�4���+a�!���J���ƓR"�m��w��C@`����F� }k�uQ�ڋF����(!!\XH��i`>o"�Pa������H|���6�2	�ִ�_RU��l,H�hP��Ϧ�#e�X1>c�}o&�Kύ=@�iq%Xd�Pyn3�l3n.��j_��%擮9W^�l���ڍ8�d�wO��a1~]�E���!�P���_�}�c��� ���~����9���g��=2�T�����/)("��>{1u��2�"�I�� �FI�8'��ٓ����8��|�:��w5٭�	>��;K��]`%���F1���[0�Q�]"���ͧ{�;$���_���1y��
��b2�L��U_�^M���7K��]��3��U����_�R0�O�!|i["�W��N�e�0��A�#�| �5�)y.��p��#i�EM���z�$��A�Th��%��f�;C��=j�yC�H`��!.�F� ��i�+�z�I�A���}�J�Vq�Z��g�t�s��f��X'�S�^�<*~�am���T�#�Z2���t���'x#i����cn}d�L2j���̋�\����!���
H�E�Ve�ERC�u���']+::D("l���ض���Cm��Z��8Z��hz��A�˰���?�/oXA�mE c��(�	g�Y���Zə�g�4K���k"~�����{�L��L!L���j����{Ѧ�EmI��|���a?zB����;q�4�����u���f������)��4���a�'M+�>^�E��Y��|O|��1n��%���\0�u�W_-t�d�a�!N~!�נP*�w���UMn�P�����q$N��%��x^�zk��\����,[ JV�1u��<S۸*���AF+,�m�;�ķ��u��{�����Xlg��!Ӄ-ɛ�МS��Y|�7F+V;�L�KJ�-�\v���s�Ie�8k{�s��.к����`�f(����R����f�_�h+�3��dp�L��gz{��Η��*)/�����Z�S��xL�~��XV�p��$x95�{�bG�Yz{m���8�#�̢�f��������8�I:��o�-�1���$oyj�n$��~�a���i��Q!@�h��A�7� �D��bX?���y��� /�
XS'�i��cRL�r���6U���e��Ԃ$�_�Ћ�Y�æh
^Z-�����&Ӿ�а�_�gy$Z)&+�/k��N7Ϛ%��)&arM��b,M��p�M+�l ��	s�#"��;],I����*Ǥi�WE�օ�E��hvʳ�������g�J9�ɱ��52gΔnWַ�D.:��?*�D�qup�)�,p��mW��.�4MK�q����������k��:�s��,���k�\����nFq����u��E�L�Ι�د�y�����;��,�h� k��ƹ�P'2�m���@�\��V.t�=s���s�w������V���y#�!K���$�M�&U�"�;!'�0%uTX����6ͺ�\q�^WqՄ�ۇ~1.Aâ�㦦Cu����`9v�tmm~���̗ePn�6j�hx_�E���b��n�z�n��t��D����ae��Jj�����<'�B7�7�{0A͉�V���b}�tǬ(�^���z��𧆔�?ݒ�W�"��ʟ����ёW�D��@ΌάFs�����Ec
ƌ(=��V����X���Ӑ#�c�������P�;��tvա�s����! ]$/��c^��6j&�%)��k�͗ ��Y���i�"���AAa��3D �oT��%7�7mlI$�6����$�d�A��D�c��͞<vޗ����Cs��U�`	.���iQY�dc�A��?Iɰl��dT}S`���x�������,���=JS!�!�%=;�}-��ߦ�1�l�AJ�yA�F�9Y	��!V1�e��1X��q$R�
����j���/�:�������4�H��%l����y���83]|j�I^,$�rh>�6Jl'��Ƀ� gHĬ2��FKV��f���iGWs}��=�d�Zx����꺑�B8����S��(�e~�D��]�l3����ݟ�e�v�̂���rF&����'�g����B4ba�$\ٮ�6�B,ԋMT����PQ"_�Adt�{�xr���Y���A@�����b�i>����+�����r�)W�怳�t��	��jx�y�h^��\��$�_���38Vl�0�V}@Z����/ 8Tȵ>c���yG�SU�kd�EAC��
E" }�����&;�3�7f@$����'��Å�N�w���M�B�ƠTy��r@���"+�4"[_ĂIC,���L�]��2�I��h�&�@R�Tצ���R������������ͼr�^��q-��\BH�I��겖��E�*���8bw����0d+n-K`=���ƛMbM��j�p�~'�~�c��}�����IW�	�"X6 9jC��P �ڷo�B��u��`y�!�B �qZ��X_l�΁x}���6��*fF��mö~���wH^Sc�0kcZ�ׁ?]�'�OV�hI=��pϰXP����رɷ`+w���ڳ���ݰN+{�Ds��\��� ?���,Q��H�K�%	4$��'/���?���dZ���[U���+ּI�p��|�Q�R�49�ș9��n�<�V`���I�a��&�y�Cq��|���7t|�-�Ef��ĳ��^L��H�U�;�J��w��O��/һ=X����ȩ��p-p���~��y����1�EO��1�f\�H�F��v���i��"��W���O��b MW�����*om�[0iݮ����R
�}��d	��v ^��0+
`�m���cRuD��h����!�i`��d�	�{@��8�G�k��[�l\�Lp�7F?z/�w�%�z��	����y�O]$�0��<Nke2��ȣ��(��o�7�/ T]6E�۔��z�p�1@�a�;��f@/)>;#��!��6Y�V�A�וȹ�=Z����a���3uM1��O��������j�_�gj�+��~�2\E�"��.�r�#M�'�z���.)F��!������2�D'���M�6E��[�J�U+�bU�{/����#��M,�~Ѵ0&��^ϔ�C��0c'	��N>����
a��9)1;��>r�[���5�p����i�@�a�(t��V�ǟ�Ц�-�_+�F;�&G�N6���µy_�F�L�Df�؋����i{!������5�V�}��d� �L�-Z �|�}3h|�+Ƈ�/��1�Jka}�a���Kj�y��9j�&.�	Q�R6Y�M��BǾ	�;:�F�x��>/K�KW+����W��xq�_��dR�mb!��r}��k����A�`3�՟�0l��$r	?���w7���sxe
kr}E���������2Dj����
=��K�p�'�~�;�lK)w-��&ƒ}%)��ᾡe�v1X2�C��U�ݬc:�	N�*Er64���vp�uX�E0���y-D5At�f0Q����!�8[��*�������-b���5��Q�g�!�V[쬢D4}�jǦy��\��'�(MT�~
Ǻ��ݴ�M,����8φ�k�v�������1W�|��4��h��dfv�/�a�:�l�2�����lT��k����.�Cx����j^��0ͺP�n��P�Zo����A�~����'��G�:uMu�G� ���!�X�n��S-��Z�!>ݞ=�y�Sy��&�HWm��8j�<wBl�G�_�?�i�������=��g���O�  ю���:	R��eZ^��i6*Ғ� ��1Y݄{�G�%Z-�C��#�z�R�T8�B�֐r$%�\_8��_ҕ�l�Z����
��!-�1\R�<X��|���K�Ĵ��0�u��@�����eM�ĺ����0I4`��.˻�ᤣ�0p�r����^d��䃑�pA2O�s��>3S&`g�<s�~�u}3<��[��E���8"����?R$��S�r��O�̋!\J4<��A��� �ok̄ �<yD���1�F�� F,gM���Z��D? ؆5��r�ӧ��AT+�>�4Y���q��F<�Mܸ��j��K�&�_�7��ޥ�N��M�z?��B���d)�)�A����#�x����j��S�;�y��]�/0�1���:]2M=*��R����̦i�'�e5p��s$F0�`V��7>�qɻ5m15�:
�+�ٔV�OKR����"%��,2�U�]����E'��^��uVG:Oa���#^�5-��5��y�a�TΉ�C|ՙ�6����������soxR�'^*v�V�ԤZa�n�%`�̞7.'�\.OuHE*�gu]�Y~G3![��2���.$5l��U���"Y�X!A-��x�9B��$׸���T�E�ӥ�R�{k�\/�E4XW�|F�e��'vS))���ɂM=R�W#a�0��=�5L?��l3e8߸���������3\�(�׷��-������6S�����VF��\,Ӻ�~���F:�0Y֥���l��2�\�:F��J������'��_�������J!�2��r�B�)�1��w����z�sl�'|1��L�l9��T$Feܤ����Дo����Z�0S$5�څ��v�1e_���J،���R��_fk���q�?�4Dm���U�L� N�HXq��z�T���N��K�A�)p,>?zy��o�l�ܢI���ĳ�e����OO�}�,���H�Y^���Oq~:pik[�6�^���h�b/����&d9c�޼um��]�~Cg!mdP*�ƛ�΃/4�X&��FN�������DO}3���H�b��۫���^c%]Y|�a�����u���m�!L�j�/ ��E&���w�8&>�a	�܄q $P��[��0���lPj�:���� ���'�IR����r��\���A,�_����ɪ�����۠ϽK�|�l��I'�:V'�'33G	���$s���`'�N�X�p��n�tݖ���ry��_RI޽�`������X�ʽ������:x#0ג�^gUE������/��Df�:&&�_Gn# F�����-�\�Px�����Y�������
H9):)
�b�p�d��ωy>~2�W���{Lm�aA�6S4/k���&�ߑ.z�ǉ$���!�0���v*��7�������8�;��Ev$��n��n�|��ӼH���>1��V�%)�%�8�S�A�U�l��:"���T�|�Ԫ�<6�~�C��f㟆���mY1E��m�
��feW(^- ��S�)rf�m�e��e�QLs YQ2N2�B9�ۻ6��UX����V�%��8���X��U��B?cugD�ӻ�2���p�m�;���2r1��\}J��v���k%>j���:�f�S=�N!Wz��<�p���b�;=�����TG�ׅ(��Du�E�"Ӆ����T���y�m���l��_A1"�^���(6v�F�M��ʺP��s��^���"* �Gق�	NZ뤵'�S˸���G#�r�¯��.�4uJ��N�6cnM)�9�R�9T���$�I�a9;��5Bq<=�^:c�3;@Ǳ��0-~ɰg�E�-؜�C�}�\�e�<���V�o�tH=���$��˪�bj�s�����i&�b.�
���2!�1#�|���A�V��0]uZb���~�����'�D�_����z��]-cn�~�	�)�|B�K(4%qq|�fF6��
��\ř�^��&g�[�+
�!ΨP��@�}�t�0u$��BW�}�ѿ����8ID�g:���fl�$�tj�a�߲	p%~�o�x�A�hy�IT@����lrFv�_�,��s���goeۤ�;�zЏ��i�+�rڊ�:�����|{7��+{���.�ֆ�
��q����2��~�-\�{ڪض��M���SR��Wle�i(�6���ןXlJ�k�ܾ
���R��]�L��g���%c
h�n�҂�y�*CMmP+A3C��!+(�����/0�k��Y�����̛hj��VI�hJ��=�c?����TgP���צx�5��s��7<�4�XLi
yR8\B�����<�Ռ8B���Kʰ��r����m��;k��x�Q��c�ޑQdd9��ʎoC*��<��M-��{\|�A��I;��pʽ�H)���[��cn^{����I�g�MdPV�%�`��!�"�:2�b�,�%q._\�~�#]���cFI�u<��L�be��k!
��ȹg�.w�81T��8�_|R5�מ�q12�x����N%�}>�Y�e�l3�׋�JP��g��)x�n��18O	/�J%�Gwc�}6i�:�Ŷt1���z׋˘ra�{�=�C�����8��8bk�ˋ�-!GZ��G]*�i�P�b.$]������bZt1��=��f����V�%��5_$�D�!�[�y�}��*�H\Ā��ɴqЧ���>Ob_u��H�z�&� i���I~BĄנ`�;��K�I�ѻ}~��/�E���[����\r�A'�P����s�T�w(y"}�&��+�uI����i�K�}��ҡ�W�i�O���ѷ�J��b��8'Q��Ƚq�U�
�v̽1u�@�:v�.E��u���4Ĳ�e���MrM^B �����MU������!yd��M�]���bG"MF�����g(�$��\�-�4n��!%�Ԛ(���l��;�	թ7~�C���	��#�dU�Tެ��٭�R0�(�դ�E=U|�8���Ђ� T��A�
t]���� ���Y~�7 8烠(s3V������qM�^���h�3@[ߎw�d�rc���f�?�zM���U*_`�`�[��e^�,Ġ^��!��R	�p�R�n"敊8�JQ��z�f�S��q3s�F�c{��]��'xM�h����V��� ���ǖ!އ�(��:r 6��ռ�艒'.�I�f�S�ev�����`/�O�����}\�.Hu�jA�f-|�!�m��Z�x�	�Zɗ�R!������]���
~��Q��X!�+�׈6�������"��V�B��:6o���
u������mlM��A?�\���tݻ��:ا���}����z����0T���s��ﰏV�R�����V A�����SM��BH���Q�xM�q#�����y���[~%mȭ��s��HG��4����G�u2u�?�S�9ᵏ�H�(��ǝ�z�������|�X��q���� �U>�O����DM�)½8�w�nʮQ6�+�F�ĞGb|L��H��U��w��疗�G%�|TbҤ�Da������i͏;xc��̸�����So�q�q��Sda�X��aX܅�.á��̣ӑMַE(�$���ը6�&pY��iPA��Y������3��;w���Q~ 癴|7Kfv��lD���$��3��;w���/ii�u����5<Ґ�ɏrT��L�yw���
.��+�e�኎Ĝ�����h1A]���x�U�iU�����l!��H�;K&�6�� ���,�h�w�O0y�<y���VP�yY+��O��9�G�/�-���P~Z�ͦ`4L�d�vVqƖ�ѻg�Ee/��Of��@P�`�b�m4�k#�i��[��ǭƩ��뾳@e:+ �%��z߯}>U/�~�#x��~A�:�����>N��5ƴ�-b��>���8\P�B�|�4�y����Y<j;�&R����|ϨjP�.na�\U��PQ�Sk��ӳXͨ�V��D�6rD�h���j�Z���a� �X�P|�~]��nv�.�+�z=��L]�|5�������&���g�o,"3�2\j��3��t���Sj���<b��>��]_J0GC2�@WC6��]�����a}��܄'��k=����C��w����:�g�~H�e����N�*v���G3�i�4S��̂��>����⚰I1 �Y��)�=�{1�Z���&̦�@v�׈.:}���U.3���@���ޤ{�Ż�\	����#qȲ˕���9�wf���Q��v�1��;9��e�-r%���ܝ����x B��}��4�)V9C�W>�`W���e��+��y�<��9�l=�1NYY��u��ˢ�6�`Y"ص�`3O�HR$�,-o:f����@�e)a���$-z�-���>�D����%�Z�5?#���2���˜wm�$H�TK�����O{Ԯ��3_�	��B�j&&��8�娅�s��b�07U�d*�f��6@~+"+$��ϣ�^3���#^JN��)�Z���-os� z�AS��#0��׫)p�z#2y�Ůf����Sz'�� �]`7�F�˝X&6Nk�$�}ͿF�e��T�œA�n�d����?��`�0�KJM��̙�Q\�5�E�����,���:%�|I%h��h �B-k�w	+��>���)Wn��{H��+�o_溢�a"�2����ѥ|O�b'�^
f��5*��	gi�d髍Si�!I�ˠ� ������Zk�q`���Q��8A����v�L �#:�5Ŝ��(gS�8��_</���Y)���gW`!�ze�e�X	VO"h�1T�{U~b~�;�s�j�n�F%�?������`�5�^�.o��|���5'e]������yg��B�O�ì�FXM� [!���^ａ�z
�b�z�R =";K
��=D����Nct���C��H�PC��-*��Y��]�KT�뮙�5�p�.����c�>�׉O����������6ء,�V��~b�j���3�72@���t�O�=����F�Ns�ɺ?��l�~�<us=`SF�v���Lą� ��59"��"�k��K."h�%j��(��'�v���J\��f��{��K�V�"�};ŠoV= �+�I� %�op�xv�`ݭ����bi.M z��^Gj �ɖ3����^ߤ���G>�#
����t1��>��5g����6��5��B0[��
;#18�C�Ð�BԬ�]���r�0�����M��>��6a�3ck>��j���Z�d�>jϼ����nW�tLwXc�D��Fp��z����cڕ���$i�ҫHz]d�����w�6��gU)x�P�I�d����S{J�������H/�ߌ��O�Od{������1�-���G��ߛ��y�췛ǯ�ʶ��>r�MV�j��ł�V2�-V���o�IOk��������=7)�}�Y���e�N��#q�HH�BK$�Uu��A�?l|�)H���:sz��ʮ��K�tcK�)���Fa�+[K���)i*�iF"G��_[�(�׵Kk�	M�� ������O)�ë��Ct�ܪh/�����S7Od3�)���PO4��"�H��Ũ��X�j��M�川��Z6���t�%4�~��)�h������*r�Ҩ�{���T�����I�]#!����;�!A}�;��v/?���܆��M����ʰjxFT������Eh�ʹ�����2��g@w�,�P1�Җ��S�]����i�\Nq
_�;�C�B��ٙY^ޑ*:���,�� q�� ����7n0N�I�f�;
*@5^,m�:!r�\-����nEj��S�wo�X��O��W���`o(���"��/��i끐rĽW�ƨ����̎�\�:�B�'
���FFaR��m=R�4CG�Wp�$�e8"������/�ę��H�k��Z�K���2�_M?&���t�0Pr�ifQ�B��]�V��,���=d�^!���s��3��o��)�]:{-bNs6c9��^U^Iʞ�Z$�V��� l9�����#�l1r�mz���?�T�/�ϥ>�z���=����u��Q
Nq^B��G�`t2�����L=�2q w��%��9+�Ԭo��~l��9g�3`T���+��w����׸�������^�88��:�ވX5�Y��)��<��`�L'#��ZX��p0Rh���B����}w[E�=��x�Y� �V[��HZ\)s9���0#B9&�L의�1iMH�\���9�ZF�^C��y��b ��x;y&حλZKj�e~� G"�y�5U��)ܦ�9�4-B�4AlHk+'���p8�b>��Z:���db�PS|�[Մ]�B؜�Sx

�n)�����3*C��c�x��7@U�W儦$�x8Q|BmC~Jܼ���=T���%h�,Uq��#:b
�*"#�Vh�\!�����'2��oXmZ�F���S�4 ��xϝ$H�F^[�cS��*?�[�".ؽ!o� �����oI�	�,	�WD�2$U���+Au�ҋN"TB���B%�v������#/��	��3t�r���6�=P*'�в�Gx�K�S�Բ��-��!H�+ �Z���@�~[p��mn9��-M'c\,gs;��V���l�{���y����D���X��h%��6��HZ�,Zm�V�ɞ�R���!�;�N���#P
.������=��/��C�?\pC��'G��P� ��G7��X%t`�{'k��I~N�e]{~K@"��t�(�CEK��,�#|�Ne�$1� �r\�Ld�C/5h
ZF�}���p4����w��N�НP���F�$3c�w;yZ�Z��#&��?����,�� Z���Лl%5Do*��:�0�@�4!�%b\F���o� T��&3~t�����j�IM���e��m���҆Z	d���K����mF-�oPc�>��Y�?F����F����g�%��$tw����(��
�o��x�m�Ϋuxp�P�c-7E�p���7��rO�	O�DE�� �qp@��2����%$��(fg}��C��M�@�gS��~r
)�:�U���=ɝ`5�:��t�Rr���8y�Kr��dܽwL��l&�|CK�Qt��A�)��c.жc1�t��Ș�c�Z6�:��5=�2G�}����~&��Y s���5�k�Avl_8�c�{Q�o��	���Ϗsb��=�p���qЦ��-��_*]o�����6	�w�M�$�_��&����^�@�����ɷ�>� :��9P[��{�Q�lW�k����n<zԮ�̘�1Ɂ��}�D�
�7<&�0xG�|����y�n).������ah�w����q�n�[�Zfk�!�,�0��{�����:��+�������Pjں�:Ȍ��J#\0l��O[���YJ+�DqqF��
S�Ta�7��)�~kQ�9��)��p1/�"�H�(�:� 󸎨�Dz.��yۑ��1�yh�i�gJ~�V���f=�,i9�ȿ�Q�K�J�*��1�}��f�Ó[`�@��ex宝���,�$Z�ޭ�^D+٪>����,7���	����AJrG�S��u�?�}�����m���G�Q��B�/K6�:y�-}B+�����ʂZ
S}��P��w��ꌮJ�1�M�
�|l��j�I����d�*�IEFT�SYX���m�DwL�)U ���`��%g� ������ބB�5���*�ﯷ��5�40�2���iɲRG(	n���i5 �����	>�RPݕ���-c��l��q��m��F�0]9����\�u�����P0�7�&VQ>��Lv���B�d�&��Qu�tz�#b��"�sŀǭ���D��T0v�~�>��������%i��uZ��՜U�5��aq�O�+��ڍ�O��1%LMQ,d�w�E��WT�	_�w��!~���cR?����tڭ�������d�?�*z}3Z;Rc�����5�t��ܐq'�4? |dD�씾���s�P8#t�h/���9���"K�������L����*㈌��3ܥ?�y:�f%�Ԕu~�Z�vIDŔkL���Ow�e��n�Ӡ�'��b��\����u�f٬e{��7�Q�k�\7��)��GR��
��ѿ.������)y��[� Ԯ�3x�:��Jo4l^���:�`�� ���'j+�d��)��ZD�6ux�Ap���-"4?��ZM�+|��6�����u��P����-��>�F��S����$m-
n�TA�q�]��G|��J��Ek�i�'h��'ڗ2�!-��2+�8՘z����O� �|�� �L��qw���=C�e���F�Q��4�+���=�Sx�X0�A.�ő�V�"���Ġ1�<��(�#��UR1�M�UM~�eհ#	l�޸��;ϛ�Ĥ��������_b2W9+I���ҽ�,�W��#t������K���h�`��D����o���^a$�'x�F�J>���sdޯ%xcI���۬Τ����8,�y�U���@d��`��6
���I�+���3�Єa�&т=��⊡��I�&�x��3��w�9��P
ur�	�ζ����'�0�� H�N�V�~waN�5F\�7(h��P�Ph����K�%�P�$�e�f�8K?�a�S��SB9^��W���x~V#���K��2�jP�o���e�{���H�k�'P�n}��ƚO�MpR���b<�>������oQ�ؚv�"q�.���+��ն���"�
X��A��B��@K�7*(yЙy2��^0��H�"hf�QQ�@S�v��fL�g)m���C�%ө#IId�^����~LusZ@SEuKYWs��go?w�?:�g�Qۏ����^ϨKܧ& t��
v�m��cW>Ǌ�
���������		$G�x�D�]�X���V��=K�w葒���)��ϘP�E����Թ/�9�Y�K��K�n<�Hh����ՂT�����D�*[
 V�~�4}rŇeEu�JK�����L=;o��6��Cs�zm�#���9����^�s��}A݃m���͍����<���[��K0���٪����׏�� �ޭ�T�"k��`�o��O�n
.lh��S".�����l#?~�����ROy��j�3֪^�� ܖ·潢����N,'K8�g�*˒�n����4��(�xӘ��A4�x����?!�q�IS�8t�=Z;ԙ�OY�0�.���g�XU��=z�|B�����@Q[۽h���z,��ج`g9
;C�ڥ\��E��b���E����;U#�x�g!,�W�I��]{?(���76^�h���PL*�[��R�������3�{o��g�m"��BW>"�Ke�� T�ө��T�8�*,��GN���`��d&�������d�>og���ϔ�kS��#@e�:h#��w��̝��C��g��\¨��E�B¸`��f�4�ʊs��[i|����mH�v!k��;j����	9���l��@��:���u����-��!2��U��=�@�p��ar��frk��h�0Ϥ�
M9�E�s��:n5I���~��p��V
���S��5��n�ke��G�	Џ*^t���2+~e�&����֋O3N��O�Zϟ$�h� }���&4h�8�kA�$�g=����-߄������M������۹�Z����>�o�?֘g}���
�zp$�3 ��҃�q@�D��~.`"�����ZI�	�nю�3�˥X�n��R�!m[�Z�;�k�j�����G��\�`'��3�l*5$�_� #C�������CT���0mKo�TAx��:&f��.Oo����p�X���j�^C&T����$$��b��;I˒�GZp�!W�yL��G�6����.�y۹��-M\��
xY�U�'9R��ږ݁�D2����l�y��:�Z�5a]lQ��	��+��!��c�!~N��qa�{Cy}�y�6���:���YG����萁�\��������¤�����uL�'��*L��^�uv�G�3��n����}s��txɒA	9��ޖ�9���j�W���k� �ճ+��0�UCAe?��Pj����H��|PK��G�H۷7����~��a�uq�Ì�G�E
s���F��H�jL�u���m~(C87
�,$��B�*� x�J���r�i���:��r`d���{�K�P��p��?�=o&�nV*35��NgYN�X=5�P��{
��E�c�&8����J�x�l��C�9F�{+�	ں &����=��t��H�Q��n�#��S��/+bـ̷�g��Y�u���$�5���"k�ʅK*�T�
�?@J�<��D`uZ��a�_�(w��#���K��.�u�GZz[N�Q+�������ϣ��@26S���n�x��S���K�����(��%�����TC��E�II��"k��|��ӈ��Z�]�'�Q��8U�$��u6(��e���¨PЀ��!�wG�&�f������a)ኻ��+'��-�TJ�<�\�C@�y�q2�?H�*Ъ���k��c8�Xѐ�|�ťB�l�AC�T��ݿn<$����������d������/䞇���K�>�x��'��r�ָ����w��%�� ��+�)mz������Xf�����(>�4G��eӼ�BN���b���OsWu��$m-���~j�B�u��A{uWwR��Ǝ�ߧ���o����K�_��e�O�l�7�t�<3�lO/�D�������bkΑf��F�26�b�<T.�h1��/�6�h|V�5�@�4�{�V�⟖D�!;�=@|���u��vA�JI��
$+�p��Z/��$Հ�<������6��n::�c6=��v�x0<��܇3������z�$����v�Z7���	�$K�
�=i�턁��- ����5]&�VZ�-��Z�	o�3�<��'n���]��k��Z�ǩ<���R^B @�)��E�d�Y'��r�'@�Oeh%Lچ���1ҳd�`���H���ncxyy�yuN����l��c%��a�l�Ho�&3vZ��#�lҐ���%�����aH�	�l��/<"�	����t�A��"-�~ǰ��-�F�m9|#��;�r�Q�ܝ����ZE��o����1%�	w� �wdZP|gŕ��AfQv�Th����RUC����l�
E�%-<"��z��ʏ��J��t��*:�'���]���͞�UMv�:%�8��_�&x\m����,`PJ��H�;s)L���a������@�x��ȯ|d,f�k�GˬL����z`ѵ�)4���f���iU��ڽfE�"8"�-�چ�;ȣ����1���q+����9:��@0���������z_'j���z�7�>�A1�m��C������M	��:lA)�b6@����8�	��Ȥ�\�U��hc2�X�c�5�Z�1�xA;T������oc��e�N�����5�j��x�-����@�
��U�,	Y��۠����fՙ�"����b�t�e�2���0�n<G�`����j/,��B�H/���~��L�m8��$�a"��%�|\n8����?jt�]�8掓K��h���#ӻ�o$f�lTv���ܵ��@�x�NZʥ *�0�ԁ��}�F�s,�\|p*��OC�I��WL��&����(����|�)z�}U,��!cOzx��"�o0��|m%����#Иz���p��&f'�Sd�� ������7���=��iל=�~՘�1���H�|#Y��a�,�h��W�)fF����ٳ#�.R2lz.�,*Q�|�A<��dؖ$Wo���Q�Ha�����n1�|�-���U��pm^��8�=����yv���kv��^��+�;��y�M��
"���mN���S��*�)m��щpEN�m+��h��j7f,�ὢ.�T����[�yqd�n��QF߱����Jrl&��*�-��a�f�g�4E	���9��[�,K�������;:?����� H���com�ô�[R��^;H����i-�(��b�4p���Ѻ61a�;�z�$S��'W�ѿq0G�7$�����פ�~C)������y6�Z�߲��m	ـZ��|$}?S�<m5�T=�kF8�b?x��Q3b>��D
��3$8�+Y+��[����P������&������1e/	c�ߩ83c�<HT�+���ƍ� (�[�|��O��=Σ���_~Y�B^n�0�y��G	r|�%�Ç�ԕ��gQ�ۍ���Ē k�[	�J�.��v���a)��& %M��z�Z�0��Xv��}}�~n�.^���-Q�������W<Ub��O���b�Dm�	=�qOs:�k6#tT�R<{�`F2Y	�:���А$y�ҧ�!���6b>�1���(b<L���K��Ӆ�''I�\��@Ǧ�3�u��o��t��C}G��-VY���.��.JG����*")�����݉��$���-ԉb��ִ�TH�Zf�f{��Ss  )�����5{�1����R���QZ�ʓ~����5��v�,��e��9G���R�d����]���=�0wm��x�;?t����5ϻ�|�w����4M_�0(/F�e����ۼ�j�u*���}����;�&6b����=26p��Hմ�]����u"b��4�
��;AA'��&od����[�7<�?MV�,����/J��mH�~��+J��)�1O~w��t�3��Ƌh ���4xja[�Zm|JApk���;�B�Գ��٠r��՟�򶭡O�B��g�����صF�����v�a��?��V;�)��C����\�1r�#���$�r�[�� ���L3���
�zOQUdY��m��qo`o*E�,.��` {���}Kǖ� d��b���@�d��Wˌ�6l�����r|�E[��X�B����b�^F_�4֡?S<S��lI.]�f�hU\nkˣ�E�G�$�ǲ�����n�Tb,%��y���e�T}_	�ʠ�H��	���]s
�잺u!vX��H�9�xA˺/c��!4I�΅o����G���GbW?N>S�Tu��&t�3��b-���>ںk��9���'TgoUgS)�?��~/Fdmo!�L�	K�v��u��L�}�G �W|�h��d0��zRй�s�#z��|�pK��]��s�ӭ�ౡ[��~���`К�j���]�� �2�%X'20�eG�k9��}���Qj�(#���i
�p��SB�=�Wh1ge�U���qs�P�6'����mk�Vm�[rJ�����qUasg�j��0���ł��a6���ww��0���J��x��fJGՕ&�Օ�ws�}� �A���7q�X}�*/음���U�b�G�.O�2H�ҩOb'�8:��	�I�xZ�R�RS`m�
���J[JtJ�
d��1�q�hfl\^��
^fMc��[_�_p�N�6�#��Q��A\+s�Iʝ0LT��(�{Ч���7"dz=7�"�E��w�q��w`*$�M����X8�,^r�d��1Bb�J�l�e0zw�A�ϥ�hq0b�!� Y��m�Y�3v@���=�+(kš���Ȕ�}V4�ǉ|���H_|�r���R!ߏn�=oPruoX����o���
*��aOA�bb4C	�5plJ��K�OٮO�>�]�2�9�GB�X>���|�]!ͼp9�1���$LK�i����U�s��"!6��ۥœ�A��C��w4�e�ﲑ�������Y�����J�w��M���qj-\�l���v�k�XAA�,(��6�ZXqƗEYfI���A6y���Ϗ����ohXPB��m|&j����G�K���o�	�}��3����(A�Ȓ&7��ْ�LV��z�N��q[�h��z?O�Z�
#=���?D��*IH�,�\�B \_v ���Q����r2v�3}�7��*�y0h�t!���\�,A4@�����=�v�P��c۸�,F��P}�w�Q��=�V�=X�MV�t��{�	��k����$�p�:$GWns/�X�F��?a:��F��O��w<<�?�d$3A(��~n��B��'&ޠ�`Y��Z��&�J8���^:���x����S�*�ƕ� #�<���R��ze1�UR(Pq�n�k��t���tTS��>�kk�Z)�;���p�9�P�UL)R���aR�4Y_�fQ�ְn���x���w�Q����ǭ����ZΡ�-�5q�d�0W5��hm�'��ܳ0�̯kcb��?u��������VT�
j��a����-�7+S2��A,�����3?#�{f~SF�*��Ru�jt9��:���xT���f���a5s�ȿ���T��C�}v��S����% Ś�3>\rI�����Ƕ�6��H��С��F���):����:І �b��(N���S�j����Ҙ�U���T�W��\6'�@L��:e4I*(�z��;�y<k�����h:Ĉ	�icNuP���Bq�S��Vl�uh�Y��'� "���V��|�A0m��W]���E;�s���v��䧉m5�8Ƙ&�ou��LS�4<jӔH'�N��)4Zi�Kx���p�+�ɜ-�_�)=^�-�Y���p���z*i�
���N��
9�)��Ŗ"�$�}�b0 ��۽�W�
4��D��^����W���G����l�{�BY���ي<�]� �M�?�ef,m}+�惬��M(4�֛X��
f[
���|L�������UPy�e���MxRW�1���
�l�~M��~g��:,����n�w�@�O�<�:7�aP/x�Y���?S�H88:)�Kی�^��<Fec��?�h&�Q����c�Ԇ=�Ώ���)#M0P�hY���*CSD�x�w�~m�"4�c�K#?4�FH�y��B���8���7mr�k�}X��D;_;á/E��Ub���S���o�5�h8=Ywi�(���&n LCQ�؁%���.���K�uN �c���ZOh���m�4nʒ�KfK�/�1��`DSR����|d��H�H;��{
���4ÑO��Z0��m���w�/6����Q�Qa�g����U4�K�&s����R/ԢX�������d���+�NֳVXa���M'u���������6���ı\�ֹ���3�+����o7²����#
D����Ɣ��;�'���e$W࿚�ޜq�����w�i��E��(W�<!����*U@
�xs�j�֬T{�{�[��A�� ��u �>Rɖ	o�E�����!Z��1�� ew�[XD�I�C�q��~ש��}���+F�^��ۗ�'x��ܛ�Y��A���$���&= �a����H�M<`4��t9�-��Pb%�-1�V�#{����w�������|�m����(���&�)���2�q bEd�1�M���U�m�9�B%U�f�&*��+��, ^�Y��`)m���A�u��k��v�B	�u��{�,��Qu܏��ݸ39�@�5�k�]eQE�ފ��|p��@��B1ɤ>����	��(⯦Ć���w��(g,g��E��L�#����70����_r�
[xX����Y����?w/[$J@��H����F?��|�e�]��D���쫷���n��9��[���T~�����[&k:+�$���g�^L�d�\����R��-�%�"�c�G_�}���:�^�ܞB�f�Z�.�?������Q$xC)V�O��,�j���%�Βk��%\��c0���ƽ~s��b��)G����R��wK�?����/�Y�1�ys��ҥ��m#��at�}�� �s��B%��O�r�9].`�
��T����N�=6�9T]��'�Q���<��t��/�М���KU3�@BLi��U�۷4��7��9����RR���h�����`��C͸���$S���n�;8Q'��gf�PK�a>��	��!Ns}�bF�~J��Й�;�ߕK����[�z�6��,?�<�=���T�{@n������׼ �4�G����tX�����ͤf�_��ǑI嗜}�i^����<͎��V�>���ɰ皈lG�������.�43��-Y�|}m� ��LfȓV�`�岖�zr��p�4�hW�'a��o!
�qh����Pr�v�����p�i>(������� �� ����n`��5�۶��T8�Dx��p@�ؙB�
Q��GYO�;P8tn��4!�`^�?<��[���s;�6;l��:o��,�^]+��м� 
��#��bu�ၥ�4�oJ������ұ!$��C9q�5W��s����E`N�BT<Yr[2U����{��'(8T"�*tr��0�f|���L��+O;�`��ճ�w��S#��_*JB���]'U����T��m���#nz�M�|C����©A��a x����]D�&�!���1Ƙ6���yB=ĭ�	Η�ʷ0��nv]����-�1I��1Q���v�4,�?1D�q�wqJ�-j@ox)�ox�v�w��6�'��!���z�w�W��\[�C��TЇw�چB�	,X�,�;�d94�:ܔ�R��F��\{/��<��-��E)Da=�x���@�N�_5����>K��m|����W
�� &�nb�5,�X����R��:� �҅L��tPb�(�]������Շ[�q�y�kk�3%K�e�k<S���-Y5��K'���id����|;m(.+pC�/҈^�⹈P�o����`��}��.��`]������ԝ�$��Q�쌦D|2m��= Ch��o`��=��T��f�ek1_��K��������w�Z$$O���<<��")=ǡ`!��?��o��Ρ1���|�W��ɕ�,4���Β�s�=�H�{l�8�{�Nb�����x3)���S
^'b�D�g�i!G��zq��D���E���_����Hx-�{Ԧ�`�i���{��vX9��7g�;�/�
�Fa�[w�NF[�NuC�C�j�6saN�
t0J�;Dw�a��qe���:��t2������Ue�� ��0/�-|����kXuN���U�@0�Ӆ�|-��4�+8?@{�՛�n����s*�;
�L)����N� g�gX��Τ�2�!)� �	��	��H��T=jI �3�Ze(	�6A0���v�(�d��E���A`˞���y�>�#3U	ż�6E�Z6�i;'5
Ϫ���.y���gk'bre���l��ei��X��:���ŭ�$��kZ	�\�Ɇ�/)��^���Hx2N6"�h�7&�/���)�|���b� �S-:�N�ROP9!Z�<xP�J�Q�s#����P~Ď���1�`�΀ۜ�Q�SY�7��n�S�G��7��M�K�~�A@�#��nNj�C�,��A�םI��WJ^$�����8�e�k)93�o�v�נQ�>[:S@�]�(ST_�}I��S�@C���M��S6R1�@%x�H��uP��r�ɈAu7/n_��.�,H�ф���@B�RF��� �
C1X��8�����j_xR?����Aß��Wѓ�'�K��1���	�/蜁Ob�����}�Vj�@��������^n���`��;̗%�;"������j���l̔U�:��j�B\�-\�y;����p{E�CA�QZ��{�^������y�!�wI(�U��l���E�g�u�խ�L���b����гK;�O��Z���j�0Lf���Ď�h^x,��Dps)ې�D�v��%�#.��@�V���%< x�Nc:��\����0R��� rA}93���ܙ��i��	?����*,ӫ7��+
O��5��ð�D{�����LSn�o�'}"�E_�8��%��90���-!���5~1C���|f�%F�*3쟯��Q����XH��%
i��2mWFf]��M!��HW�2��Z��&�ínڭ���|޶����ȆޥȀ:��h/ۖ�\K�$}���܉;r��GC`�x��K�����=�G��xP�����e5��̦��O U@&��ѱ�����#	M;>?"s��7�uJL��6���ѹR��M�?�%�?��l����^�5��W_���S�x�����T��!��������V�����4O��4�&k �t���֓�T��*z����~g��v���Q��v��|�w��p��djZ�Li%a���q�M<���7�=��8���0��j�eo�\�B:k�18��(�ږf(�t��ɚ�Ϗ'lg�@3e�r\w�N�	���	t֌H�M�>�F��|���1�1h}�3�z)�bl�;҄Y�(����8R�l3���:�t�K��Ts��������2�����Ύ��_ǂ�e�1(qxmLꏷ�?�Ƙ^p �\#F���7���dS�`Ԏ��)�koy�%R6�3�:uh�'9+��҉��|���.
���oq?"�p��Ҙ�'$rGb�;*�`\!>L�MT�;���0dq�p���j�yN;��b[��J��F%.��'�S�{Tok%�Z��!����]F �"�Խ�F����F�@�(q!�;�� ������Za]s���>�ƽ�z3M鄄�5��<�C�B�ɐ��sL|qv�}�W Bi�v�RT��I�
������˹Y�����d�Gnm��J�3����h��D�
L�C ��!�F�T �\��ל�
�yA��30O��}x��P�EDe*�c�������-Î�Z�)-�AR<]�g��)����T�]lW�t�N�6؁�n��h׋����G�܃�D�B�/r��	�2��:Ӱ��m�รEF&���w��B�I}��&*Zf�y���$K�JQ�X�8�FBJ�i��E�o���º@��y��8�4d�T&k����nٮDg%��g⦤YO�ᶁ��y��l��b	�+��\4�FN��P?�3�̪r�����}����N�(<�(�j��V�`���I��|u�Ŀy;�%3�A��9B�J?H<9�ħ�/.n�X�cE�F�W4u�$݄����P3E���D��A�����N�r/"�)�+���j�>�?S^+�h�\�մ�&�[�|OG�
���MW��O����H �L�O(���:���'���J��+o�G� ��{:�G�3O2���=���g%��ӯ4�EZ�[����%�Ib����뷞�LC��Q�_��%�B��!� �:9j:Ez�lF2k��yX�W`grQ�g�k��:����8��1�@8��D�h�n3X��O ��`L�t�ۤ䠬��@��H���kM��tAH�W��C��<��Jw��_!��� �É-�L�i���;>�D�#�</
:�I��$/�zs�8h>��8些j��y�����\3�$����^����6��!i�%2�#Z�d�Ԭ>������|S��Q�ˁ텎����\���Q[��v������g;e#}����ZЯV��n�7��|a�Yr�[��w�� d���o��m���"� �/	�4�U��s�G9wz����Sm��2���l�h�?�yɑ�����PSD拰���Iݖ�%N�����xU�4��{&����t	
�Yڕ)%�8�U�3>��l�|�u�F���SX�l�.�ha�U��s��6<��>�y�b��8���M���L�sc�l�r��ɾ�(�YV���c�V/��2T#u]�S�����w�Pd!Si����2o�����zBJSF9�����О��_��D2"�&�=�EV�b$���O�P(���L1xm}B��^�* �3c&,���U.�_�j-[I#p`�m���,`��@nΊ��D�U��d����8纁�����'3�&:8��}b�;��c�s�E�L>��]��C��Ǿ� XH��0{��������1�ا�a����tp���Vz9�i�'�p�(��R��������׻� b�R��/�qGD+ڟ��Xr�!�3im���WrM��B�v?}���T���
<z��y�Ow�u4�H��Z"�\����G�9��W�#n��o�)�5�h��z�h�k�o\W�?��[c�rTc�*����.����F7���'p�t*�3e3��/7Ç�ݝ>|�U���Ý�	�M�a�#=]�@��]�?BQ9 '�9UA�\(���(,lw�h�]RhN��Xj��+��B@S]d����h��;�אt�� {�+M.�"h?F��3��t��w���3�^�H��L��j�ȓ�tK�y��jg�w� f#��d2�Q~%���ZL᠜��Ae]��bak�ߨ�B++k�j�JeD������
����I�n�,�Z�4�[}���^1<ltvG��b�W�<)V���]�J쫺k�`�U$d���@u�t�����*���lx��z7� �&/6���)��ZJ�����'�-��Q���`�Ld�{���'�g�qi*C�Ň�^�.��l�y�&pޅ�m�u��Czi���ig���]�r.��	��D~��4!��ܶ�tq��\�Qkן7�,���n�� w�И�d���������q|}�f���>R؍i'+�$GSLW3�$�	�	~�����y��6[v�н}�h�o���3��B��ɾ�<�����KnC��J��U���o���I��}�b�!w3�]�����m���c��Z��QJۆy4oʶ���E�D���Eb?G�bY���������w�(��7�Q�����C�#n� �U�X[�11e6���P����� 3Fn��˴[(�]�I�M��;���U<'�D�P��g�J4�D)�[ǡ҂��X�y�ʲH�V�L?rM�iT��I�Xd����O4q�b`b���iN$Q�?�������|f��D�MO֑����N��di�G��W�J9p�!��?hEU+��ZFӛ�\ī���/��+�Xd����2�-��4���>�ݦ�����=ͤ�R'�D�����3��T�v孹�ohR[�S��c9��_���X���9��o�>9�!3鲸o�!�g�~�����K�쿶�2����=PϾ����~#^�ޑ���%�hB֮\YU���R-&w`�n����-�) Q����pZ�n��R��Gf�_Z*W��l���4�>����l�ƛ���Ԃ ��W�s�1����_�C���L:et�Y ����f�Z5ˇ-+4H�(�=��|+ձ;Jf�o�^�Y)Rj��!鄼*�p@3�;Gu\Ұ��ۭ�k��4�k��Pp���kV|�O>�ڑ��;��A���v\���n�AK}��{��H�N��l! ���F��R����ҫ�u�iE|]��N�.m4��o
,�'/&��.�=����0z3���:#�ԉ��b�N9��fZK!�e�ZKOXYN#�UҔ�0:^֔mHU�����]��~	zv�K3� ND~��3�ˌ�GrN�����v*ubB�]�"�e�Q�g�w���G�����:v�����CSB�}Xz��|$#(|����G�q.n�V4#[��H;1L�i�h���C���c����y}��0�P�����Z<�z��0��97��c�E�.�V�1Ox�6�)rh�5�$D�6�Gˇ���A��`�Ei��q+� 6������rb/�+��I��eK�=a�G��W:�ͱ�TsNvW��o��4�����d��A���{����c�@܉��c�)�'0K*Gf��|KU�+�j��=&�lΣR����R樸/��d�����˷֓q:y��?��њ[1�K��޽�e�yH��)en�l�2K^��_��C�D���D]�p_u�_Bs�k��w������ �lX�*�.�VJtD�-���3�FI>�hC`�����OMEz"z�>���xm�*�Y�y���b>]~�����������0�V����!֗�V�O����Bi�i]�o�7O~�3(�2��c��w�`'d̀��\g�Ʋf3[/��M�@��W	��/�h��6�c������x�{$��~!~�q-1��Q�ą*P��fo���{�bH#Ěq�ş��<���\�e�t�����r:� a��T˳�Ssf�"ʃ�.�+$n}�{��Qf _N�<���uF��A^�!�;���c��1���۟5����(�Q��ǰ:
hI�.kE6Y�4X�D��0tD>���p����t��.���4oG���+��&�8�T7��Rk��x����[I��?�˔��5��z���(b���4Ӧ:�W6o��� /���-���ɰ�8�i�L@��e&i-rb�舕�EH�|���]: ��B�z F�B��?w&�+8BxZ���6Ä٩[�� :1��j3%�`5{o�����k�PfvVΊ$,Vs�|Wbr��/��No�_����y$��}L���])�cX���2�N���� :6�ή�7+yn��C��t�M}\��3��p��ގ�cx 7��_� f��j�@ƍsa峖�=�ߵN����/oB|� �+9����� �ˑ�y�B�8Ft"����2�B	
��d��TI�c��[ؼ�x؞�H��+�u�"�5��cw8?��)8��b��:��W镂��Ff�)Q,;�{im�AF���D5�E�1��и�
Ϫz=p��[xd�.��G�NTW4>��gx���R�W���K9���w�6�l>
[�^`b�2	0���@ ZX;��f�Ჯ�f@��0;�	�d����?�>ԧ�_�,��]c�H>&(s�]�3]�鷲��t�)�$��#��c�o��Gj�ū���o��=Y?EǪF"4�W�.��t8b����B~`O9d��!���F��4pR�#খz�vj�Ct�X��fZ
<�I��� �l�I�K��z<n�����˽��<K�}_6��OwP�`�e�mB&|u�'��'�®�@	 �8�~da�Oك4�d�pn�"��R1$!w����L����̻� L��)���|
�"i��PFr�?�7�=�_�k�!��D����W-�zNccV��z/�[�Q�l�5M�ڏ�����`���Ix�Q�6��}Ǖ��ʲ�#S����'������o���!�j!����swk��
-Cx�m7��<������uC�K|s��]�ayP����L��w�7���T�b4�ǀS��n}�J��S����h��;��"Я�sYD�#��d!�ɸ���1 K�g�)�M�.Ȟ�����$��Df:��-�څ��y��5A>�D"~c3�����UN�G8Oc����p���Q��M���Wk�q��~����f1Q�`vmd��ʧ3&�����Q\.��D���ˣ�~+��\��M��a�2)�X�#���<�1v6j(Z���[c�6E�Ut,7�s�cR&F�Ȯ�p3$!�c;3�j�a��Lۚ�J�����Դ��k�N�Gջ����%��O�0��� Qr �Qnq�%��o�l��1�TB�&�à�ؔ��B��L)���v�̘qf�4o��DW�$!�[���:!y�
_���:�X$v�u*U��o��Lk<�XS��'.c�L>��"��s���-�Md��{T��~c�L���Lt�GU5��#�ZMٷc�=�t���M��,��e�Q��E��w��Eux���ؖ=D������|i���#0�Zs���,Z�h���en���$�QwȻn�e�!GΠ�4���5���X�[�cg8��(@_V��Ҍ�󢈯�}1���	mˣ�`J���$�e�B�y8`Ӣ_���_R��o�Ϸ�s;G���N��n�ރl�� ��N�q��7h\o��F
��#�D�O��n�g�)�K��Om�����{���%5�N��>����{��Y�#��m��c]>�0�ór��!8 !fvha����hyU0�����s��ET蘚q���`k����� `�pA��m8�&��(�p�?�+m�R�56�!� 3bWiK��ұ�;�2�F��MM�u��R�ѽ>ʑ��ü?�D��[@�_3�#����yvk�4DeJ��X'сB#N��4��;
"�p���oC���������І��U�/ Y�l��	Q��(	�o7��B��.a����ζՂ�~��!�I�5����=U8���٩��/&S����*EЌq�t�uF͝;wR�X;��K�W7QU���_�*s�Nnk�<Yw�!TQ�$�<�ڒN{�BZ(vo{C�h��c��t`�1��_L
��m��-Y��U8 �����/����5d�G%��߻��t�����{��S���r:3w�=�ہ�
��� �!���x�9^�I�¹�Т������z�#�vZ�f�"~ҫ��[l���f��V$���b
�S Ҁ���+�^�^�"L��nM�Z�|��]�V!�P-�&Y��	���He�hD����O�M�1�����1�����\�k�@=�V"�_����4�z�M\�qx��𕸦SD�S�d7m�jY\��R�������D��,��;H���[͍jhlv��F�g�oy��s#+���+�s�x�P<��A����u! ڲ�&k{Sy���~|�������Gw����4�E��5�C�9:�j��U�y{�cP/�CX	��i�����,��)yH���ND�
���d	b�*�覮8���`So
H�Xh����z��?�x��g�Z�O�V��ם��eY�.	�e=�E�~�_�t
^��Gp��3~�F��~?�P|ix`^��t\����w[v��S)&�u��g�zzL��i��,v;�Dܲ��AtR�� �r�o�64�K^S���!������Z� ʁl l�~f�X�eةZZՃ�J���� �Ȧ9��i��3M�]�C�@�+�HQS@*�{�dMf�gp�V�5��p3�!���=۶1�o�
��M��>|��$��X�#�c+�L^��(�'�����C��3P�R��kڊ=zCZ�M� �a�m6�ҿ	��!�������.:�~�e�%/<l���L6ͦD2Vs��]]ǚ���ƛ�N�C�����d��*����׭�n�G�Ƹ5�>�C�><1~U��XVذ��*	(�K����1H�*w��+�֔��d�eR��+q�6��O+~���G]>���4�s 57!Ġ�D�zRs;��FŞ<eޡ�4�XNİ�b"���vb�ٛ,)!�Q-��E�~���3)��'�:�p�Y�m]���t!�7����V�9 ��h�!g�/aY���u�Bj��� ��0�C�}�Hl�0� �����e,��qattF����^keߩx��	�̼����J8!A\|Ǻ�,�v��/ %�#�a9E�6?�i\�(�-��m.��W�Xt�l��4�t�٦գҖ�Y�Kb1�r�aQZ���C�5�@��xC���dt��#�*�gQ�G�D��?�����O��桛w>*_̞�����/3i��ߞ��[���� ���^|��,��n1L���.��m
ˊG�bQ�b�p�E琧B.%�Ƀ\^ �6U�ƫ�\��wC�rB�@��"�S���s�_���!W`ȯR{[.�ڬ�TqvЁ(���v�Q�yο��_�w��8��R� /�5M0u��+�8"kн�}z�ob��P�-p��꒪	:N��u��xg���y$�x�4���
z(������S�2|����.��Mo��čX4T�t���������@^+SxB� ����\Z���X4���b5���ضi�XdJ�{��������G�c��L$�u�?G�#�hF	�W�n�Es��M�h���>�kqYU1��0�dx�����.�+�z0�)ݳT�e޶)����d{3��/sq8Yy�%|c���&V���.��E��5UV�3 4�g�یΛ�P�e�#C�N����$��2d4I�ΌT|�q1_��b��ŝMYh�C"�'�-RoS�
��N�|z~2𨑊2X���Q ?w�Eק�8`|Xgخe�ĕ����B$�s���� h��!\��G��� `y��}�B��� :��pe����A���2gx�G^�\~� eI���$��.�h����ן�a����kPN���e+5�nu�?�����*�ה�x+���׫�h���u��b>D��qOQ�`ejY���2P.",���	�5�:�Esgbi�xu��|���T��RK�q;ъ�k��n9ǈ��R2�Pf��ⱻ��ęn\k�7.�-���D�/�F��^7��?�K	�F�TH�XS"��T��ᥠ2ch��m����`>|Y�?A��Bd��$jО�@��jA'M�m"�O+n�z��`&�f���5�sq��\�Ȉ��|��|���uă���֏F5ނ�q�g� ��p����ă#�I#�����x�ŗS�uƫ�I���w�����u��p7�O��f��@eZ���I'�O�"@N���(������F4
6U��6B��0Fs��.�h������<77%��[���!� 8��d��;n����ޘ{֮��dPr���j�sP����"��R �H:�7������)�,�����?�'r ��Y�����N&`�k���K:�Y�9.�<C��CaynË�[�]�O[�cj��:9i����c2u���|[�����S�>�=��+���,�Ԍ�PAZ>�y�<�-,(ן��~�y�3�
�͙�����M�a�\j���Y��N,|sT� �8�#W��SQh7���G���4��s}UxI�����Rp�/c�ϱue����R�\IyoC����b^-�<3F a�.&�ܑIb_��z�d��-��-��mS;���x�4e���zv��:1���N�F���"�\?�ɜ�wSZ�?)nf��ԉ�8��1w�kz�k��̙�̡�r�$�sVr� �yN-/��BA�;�
����iEn���.���/�R�_�.��0w���OKe��Î[���|�
����)�r�=��	���1�Ah�i�,�i9��9���o�į��ԇR)jܾm�2��׍S��c�G���yz]�yxuA<z-����>��M�������'��$IU���|Ҧ�� ���\u��{/I<ӌh!��k����`�k�g�g3���A�W��CS�k�cT���'O`T����pc�B�^�@��q͵C�r7�V~-1��9Ft�:��1.��6�'�{y�������~�<jA_L�J��������c	�n`�R�<p�g����u8ss2�qc�{O>>�V��+$�������o��������|L�)�==�^D!R��)�
�w����˾(1~�����iò����{����`�Gl0��jUK�&��T��g���F?˴�M�0X�ˁ�XQ�N7��t�Aatl����ap��X<\�s|Łm{v�s�X�QKc�P;���\y*-��Ik������yy����M�ݓ�T4;��֔Y��>���%���>7T���O��×�-��%��Jљ���$ A�((�4Ɋ>��aL��\��-���=ƍ��H<k����l�K��N�d ?���G�>@<��8L�t�h�J�����S��E�^�=�ߒ믜�!*_6����`'���cq�\N��G:�H�ً4d\K��K[�O�5r.+(S�) nHPFdϦ���&�B�"�t�E6���J��ޭ\�������� HNGq����#l�
��s�ΦFu\B�Pڶ
�|�E�7eI?�u���l��K-.dT��A�Է�$>����^����ύS�Zݜ騆��I�D��C��hmN�" ���6*���_bH�<�?�6<�!Rn+c�FY�Ec}����ն���4�c�<)��Ep�td�O�CXv�:�x���s� b�:]����Wz�a�c�2%��#�%{��oA�ؽD��@�/�����r���p��Wi�!�(-(�-�\�4��#G�N]N$n�]�>�1C�~�ߑ��C�A��sU�X��Y���:".��@ݘ��A8�_>0{�j�<�xL�K$T�Sn��r^`��JjM3��g�Gݖ�x�v�	-#l�N	2Ǚ���52���<鎮Euu�����k�0f��VVbEm�f��@~�.�8���[�;o*vS�/�C}5m6�dxo�k��s�o��Q��v6^Y���Ne����;�{GEu�A=&�2R؛�	� a��"���,���68�	y�a����9%rˏ�1D@�\~�r�����d�L��#����QÜٞ�L�yU�,!���:~�d������4�&I:f��y�"	6��ڴ��Lz~h��\eM�a˃6ɸXO������Ǡ�ʯG�앵gx��N��H�@]O���l6���$�{{|�7�����qP56�V��E
�\a��&^��#�w!�H��ڔsA�-�T$�*�'6�m�W.[�%��Wԛ}qR/L� �K8������е��WL��ง���#nX-+fEw�&H�Pq|���U�/o��٤'����6��F�g��4���/�y[������G4������
|9�'���P���Ƨ9uq#�5%aE�����Q@=:l�H��~v�Ģ���63�GM�͸i���|ȼn>M�Y�NξVYB��T8�=��B�e�*w[�.�\֮�(yЫ5`"z�� �N�5Ak�	.Kn݃=9�êˡ"�&�W-�9���\��A��M	���z�s�'��ReZ�{����c���72��q>���[Ϲ�L>�'��e9lC0�p~� ������2������:ߪ(C�����I^���?��x^���� ��5��~<!h�mJ��:0Y�/�L&��X,��y���яÔn���e�-2N��lv�$�E��5�[iGr{�I)�ٷHl�� �UJ'�Δ>>û�w{u�k�{�1�,�Rżsf���A0�ɣ��W=��9�׸+���#� ��췯|$���T�D��8-%!doVR,Q����O��4�u�w�ƪ�sW��3jb���[$x5�2�`������1��ne�emR�Q�L��n��
x��L���S0�!���'�e.1�JhG�#������E �2�
oOz�5�!�me0��i ������6��毌ţ�nۙ@(�����M��I,� +� *�{)(�7p|�)A��k�G(�i����7~,Pңx�k���^�/��{T�]�<����"!�d���F���3��s*��ft�����a%����TZ�8�ͨĦJE(�Q�f�q� J�KV�2��<ٮ�Y����Z��g��B���$�ࢭ�9�׵��\�̀��_�s��Q4F�}��m 7�2��R��RfS���7��f ݂���]��]�kT�)g��ו���o?���ɠk.q�)�8�}�b������,���Ѻ�z���b�byJ�.]Y�\�l�x���H���t���(�}��A���x��%:QX�@���d�"����!��w��1�.D�� �#L�"�8�M�)|H^,j��.P�LH���]��-�l��bVpؙ��3,�l��sЁ�TwV��^�m��q;E�v��9��(qJ![��<�{�MY[d�o-OL���HF�K��К��#,Ҫ�e�x��&k<aݜH ْ�Ǟ�kYc�z�3���a�T�l4�ycpr�Ϛ2�����Vt�s��Պ�Kl1d׆+ʩ��H5mUN����tm�Ztg�M��1�x��L)
�00y�
f����\�ߎw�z%��=��]�y�Z�#����S]/m^��a<�AJ?A_� A�]8R� �j����v_E�o�[:�i�N#���o�P�k�\ �4�y�x�v�H���~}d����b�ȫ�Na?OW�} �uM�����.T��_@�|D*�Z��i>�hu`�� ��5o�ci_�o��TW,(�*(����pc�0�#��`���p�">Z��c�i
�5F��L��C'�ր0\ lO�@�l^}�9!�^�Cݏ�߆�l�$�kk��d�U[CK�������O$���G��p�hAmK"�N��>��?�t��e�|2��/�9kf��D�L
/?�H�dG#�ԑ֨"��Cf����*����wQ;��' c�f�{U#y�%��N����@�%x�>��*N�7�g����ώC!z0E��ƽ7���٥�2�_�g����ew��!�l! �ӄy�n��!�~����N-��+Y�B*	1v��g�`�D�gA���&����Ύ���V�I��3��*�C?�����g_�j�\�(V�Er$�w��n�&6u�=���r^����F�dg?f�0�՝C����!ob[)-����-&�14-�Y��祼�a�2L��5�>��q���,��WW��5�Cy�����jUܤ�WJkK)�cy��PP�v�$_B���N�^� z��I�r6�)YCuƆT��+֖V��sRZ�n�r6=��p��(!\n'�%�,YT�]Y_���lT�C9n�������5̓�vv+���,-�#vE��_f[�Hgh�e��$�|�(B�]��wp����5:��+���O T6y	%V����޻r$�t��+�%ڈ�dF-`L�Q���	�˘��l��5���|c	'�+��T�_�h�SQN��ɯNj��Xږ򦮅C���ǂzu��aK�H��ᦦ���	��\��FxK�m_��] �����[��M,D6���Q��z�n]Hڣ��w���9�ǌ�7�h�]��h�PY��.Wb��fM�٬��p���A)��
)�S��D=��x�q��"�(��%�Ń�d?�[�e�ǵ���>߷c"�������K���)l�H0��K����� [	AH��J���Rs���]:�lvF��ʃTh2;U�e�	��)��^���W?MSbJ�}5�Z��K��SrW���ڹ�SU�34�׋곽���3Jh���a��ڽ�Q���x�+T��$u�Ο�<�]��R��~w�1H��j�6�#C;y����5���������h�g#�T)��t�����!���
�{՞��e���(���ﶜt��$�s��9(��V�����!�Cӟ�:��:�����A�h<e����'u�D�3�)g�	_>,���q�3�S������9_k�"��ӈK3�G`�vj���cj���V�O'�^���x��#x;5�(�tC��O� �H���ak�\��!�FQ���Bh>�����'_<��8gջ���l���2�� �4�`RB�� R����09���T�r���薟�B �/]Q�,>�{�6\���!`NB����!Q 5���9K��it}]K�^�����p}S�HA���H��ރ���΅�+�G�
��H����^�Ӎ�9��?���V��"0\����tZF�G����$���2��2Q�s�ˑ1A3K�:�׭���e����(f��t�K�������1v���M��Z�3Ut��
0<�����IJ �(�����i��GZ�fJ�>z�3�v�/r�P��dp�w��E�nV���]+�+#Ng�%�f�+�����8�H��� !���"�h���W&ԾIP�4��;B<�m�Gø�KTd��Jq�'�?�6�X<-1�,�QY���tkE� �-�a��4�)�Î����&B���-4(8���R�F[���?c�"��19�����Q�gǿR�䄵U��O�H����5j&��+akxyT[!�Kۺ�CLAX	�g�!���6��@c�<'-v��<�<T���?D�=�>\s"d갩�s�)#��A��`�XGY�׬T��x37F�Vr҇�h��w�+m��1���U�����a!�G}J*#��$�w=�&M�oR@�_�pem�?�M�q���'���?aw<`{)���O�2�H1��t�x��� 7xY�yS"�B`78�{�WE}p�	C�t:�y\�KN�� �9�%x�i�f����(��m�6/�AU��<gh�.g�h�%��.��h���#�*�m�1�<N1]ڽN�\-Q�ג�O�1�(��H^�(�?@�Q�p�ɑ�H
�>��
ݦ�׳�[Hd��/�E�̊�`�贔��A���C���Y���U����������'JpY����|߂����ʓ�5ڹe�a�YWu�-������ZB����k\[���0�F�Ђ����e�`^�Ǚ�Q�����Ɣ1}���1f�� Z�s(���G�T��erRT��X<�V�B����8�!�A �S���_(�P!zF��Jw���x�I�-?	�J�M^��;H,ch0?�d�0v,�U��uI�W�|�ڍ�;��ӸDG�>���ȣuN�#nb�x/`X������񁻈�I<t�y|X������-�2K�7���T��|�����9���ڞ���kq���HE����H+�u�A�w��|u1��+4�!,�р��*A�V���5|�
�VhX�����.���R�kO'�2�F�U�3 �G��:�Hxސ_ .=ܜ�+N�g��z$= ���Uh(/Cj}�������~�W
��	�_��D�c��v�T�C�b<^ө�*������^��8k]{<�e��U�3�L)�s���m����!���u/��4����[9��llҰ�)lm�W�ۏ�?��X�V��JFFo��(��'V����A��(ZB�i|KL�`x���[��r�.l/B�J�<h���ԚMX���BU��p
��I�{a�V�j�hU�'�^�7����١B	�4���5�4�-�c�}��LhR�����Ru^C����RJ����N��#�(�IȈ���􎛻VI��SG����Ѷ<���2�b�c�� ����f���g���O�j�&��*e9C�T��A���.G���� X�^%
�l�&R�-��&e����Dׅ`�)���Ң����٠]�@�Z��#����:*�PB�ki�$�b;��!Y�WLd�9l���A���:ǈ�q{�\2@�ȶ�!Z����\�W҂�����޹%�N$+��<EBD
���^M�m}ç��Uo4HИ��A[Ô�?��T#�}��1�g�%~F��d�VI�Њ�� �����V�e�2ۨlEv�߫�;�� �D>��O?��̀��"X$Q .򠻰b3�My2&ެ!\MC����y*ဵ�c�}��e�'�ޖ)�u��*?I�tz:K#�V��xt4�,6�6�W%0�'-Ϳ3�Ϯ����sg��M N�W4��9aXH`N�^�.M�c��U�M���[g�A������E@�$�"mh$�u��(JΨ��W�6p��Q�4�:1���Gg�g��M��ZRkܰ#�s�����i�0FMʅ�KA�:������fK+�����*A~�(=N�_z�
[��1���q��c��۳�2dO������t2�JO�' ~��#dw�Y���^��P%LANQ�H^��Y�/}��(�� �*�}��z�[�KkB#T��I���*a�TM~�1x����=�(pw�x��������.4�-�v��s �Lm���k��D���l�d��k����g���*�q�||�e�&��W����D�cb�#[��ǲ9_�y���dC4|�ZQ�Ě֔���i�E���e�.	nf�=�y�aPh��Z0��c^�T'hH�3���e���"�����@�ϡ�yJ����G�%�V���A�d��ջĬe��僋�VZ�2����fn���s��7������p�4_T�6d�Yӥ������{�SX��R{>e F\;��zR%�EYO'q�:fzw[Y�l׃�(\�zLܓ�.�)��4��*�F��8Jв�}ɨ���Aye��Js�&o3�u$�N�y� ���xlq����ǦD�?�H��&��y����9�K���(Ѐ���\�1!�<�Ĩ>O�}�X*�oR��9����O�Q��b'�	GPч0� ,�g O�˟߁��.0N&�k́w?:Z�`���Z�K�K�\��V ��^�Z���:�:��!�A��GuzS�d�������r!�6i�Xj+�U�Q�ȷ,B���ݒ��ȸr����Н#�Ҝ9џ��ܰaC���'sh'1�[c ��t�ⱦ�����+u�/�}V=;�7��wZL�N�X��3���c��*��e� �RG��Э)�j�jP�����c;��Q����gq��I�6+�p���e�w.�L���/=#���E���Y�t}�3C�y�3L�� Y.�ٻW�a�n�H�f��=���0lVΏ�$��!T��q�sG"|�DƜ.��,hUS�%�W���V�`;}4���\D����O�Q�*]�T ��0�R�+&<3 �#�h��>MZ�;A���ii�śݶ?��b=�}��#���2�Y���+�?����q�'�l���3�G~8P��Țe�G�N[O�I�%��zzM�̷��x#^���J�r$�4��R��d���01��>ZL��+���c����+��9�b0�P���A|1�1������=e$7槮�EX���'��p:����}^)@`��F�{�zqV�kx*��� N���%������������g7�PE�������74��5Y!~�$�^��{I|�r=D��0Wm@�Gs<������K�p����I�!�b���bkx8
�9pא�����7�����'��^�.�*��ҰU���w/��\��	�j����6x��!�Āμ�?>C���
0��{9i��F= :�`���j=��5��+6s�˒�#�����&0*���6� eUs'l�Pb^�> �%�#�:���G���K04�$�0Z8���z&�P��YT��I��4a�<iD���~��K�n��U��qQ4p��Evr��*�a�G�Z^��_�w�Q/ k�Ek����bR������ً�ʡ��B��Q�,�&�ԍ/�aꈅ]f��L�Vz�Z�^�"l�@�����w�/�^e��2!�u��YݩC���s�������uȓ
�m6.��T(b�;Y"�9g}q
�/�1f�i8vi=k	��}�K��i� ���WD�.I?<�������*pI�h����ȍ��FQ�� #��R)3^�ϖ�`g����yim���
S�È�ܧ���U�HJ��a��D��.LE������<8�ԡ$�n%3�{}�u����G�T�؍�	���u��u�Ӊ��)
 �+�W>0�����~.I���Z�gŐ����S-%��N �ZL��t=M�)L����ҊF��+�MzbC0$d9�F���I�mql�;���^RYl�ǖ¶��=���X�V>� GA��Gn��v��vÃm'qJ	����1���>@���M���4=R����.� ]E^�߉\8fF@̌�[sׁ_�n3��J&\8�N̄���c�x�j����L3�LD%@�~��2O��h�f�D0���("x�<J'�P"l#�β�j����L�ѱ�=�~�L&s�͵E���9cP�o|���̍k�)C?���F+�h�+�@���j�e/���]P�R�����޵�����΁t�7%�Z���x�s�d����&�����M�al����Iw F�Sv�NU�ީ�z�ѩ�����N��%��QCy��f<�`R�:��*I:?<Y��N��K��~��N�I$�'k�eG�.�����#;���bx�TC�9{���ԯ��A*���������#��M�$�W�,1]WxN8�����.1�,�rN�q
�4���e���30݀oY�z�����j�Gs�zd����P�NL_*�z�ľ��׶��S�BJXG��T���>��DM���의k(dm۟\4fƕKwE�B��0�<v��Um��2��vm@�fCWW��NY҈�ð�caX�;�5�Hj6Sq�<X�H���3����äR  }|�?���3G�\B�l�LL���EL��<iy��Q�	GF���Jk����ش��a���H���\>�+2p �¦����A&�9�����Ige��\cWn���F���[?�yA��B_�OӾ�����3W���~l��ص���F�rZ�ɏV�\bCW�ͯGg��e��)��ė`���i���#�KlE ],�5�S��q����8A�,E.�0�x��#{3u�IF$�'��xb��-�r\ֿxZ�(�lĜ�3�#e�"�I>ޱ�Jv��}��� -;�.�{�4��~œ�%�2�/
��Di�T�������&�XP y��簩3�sϣ�C�����]�B�3�2�>��Z�����sM�F#{G��	�O��Y���IS�R܅�S鴒h��uD��%a0�7/�	Rįzi�j��ދH�Y�6�Ul1x|ݹx:̡���oR;��'���\&�op],�MHy0�_ܡ��P�	�أǔ�&Ȩv��q�R�l V������D�N���nOu(�3�-��)Ŝ�Ju���o�kh�=��=/�`7s��*N�[�tz%�=�ЦI�k��w�)T�<��嵪�	�)��M��%7�Y��/������?�ﭱr��K녦����~n�Pkc�v"�o����2ɾ��:&��^��dF�Q{'05��T0A@Ül6��ݼ9�,Hk�����)uC��ɠѭ�n���s-��ԍ�:�9xɄ��.�#�I(���80Ӻ�r̴�½�i�ad���B9>�LI[��,���"R�$WG��9'��M\�_1��Qy�̿��ki2\������5
z:`��s��J�(P濟iQ���о���.D�t�Ø�v������W��:������Dh��s�p͹14� ���*y.q�L^�S���4 fi�"XO��X���.�e&k�s��Ry��m/(��4t�8ƀ�JE���W*�x�\ֵ��v���0
� ;�Y��?wU�##O��u�: PU�.MZu����ߗ̆���Y���w�I���d�|0t���Ĺ8��	my�L�i�@��	�gQ�f��L��c
w�����(^����JsA�H�Q:6�(��	Ϳi���!;�W���K���P��KRH��X�Y:\ ��v���(�!�(c�VO�A�ƌ8g{P��	} A9�����1��� W�w)����d��ΰ�*�e��
�܉ƂZ{�����(ޕ��Dv����	�U���U�i�问�R�ߑ�"-����*�i<�g��� �/�A^�I=]U'n����zA�Ą�q�@�!RC��t	5O~
:�Br�):c�7�,Q	��sRZ�j=��uӥK��tU6��9�'�*L���֚��ݎC���m�m����X�X@]���M��I��I,���|re|�
�٭�H0mџ��夒��y�ǆ��J�����e��x��j�յp������H
��n9�WG����/ Rd�i��N�- ;J�9���֖Z �M A���M��%	��PѬzv�*��o��ҍQt\L[���E�t���͛������{*�	`!�b�y2.�Ų�u�@gF�X(���-���>������_��la��2�8�Z�M
�W�{�u��(|����	e�>H�1��.xP����WǖŠ�Z��I����>���'�,�L���Yd�������Bl�W�v/��_��h ��/�
�`#<��apX�^ߓ m �!_śg��1���y��ƭ�:Gb1�:���a���h���@BVN>�SD7��clTM���G
��~9�!Ė��3��Ƹ�z�e�����s:j�C�JH���)����(8��e_�2���3��=��m���r7ř�@qj4��4b�����D&��"��ȫW��G�P�@5�� �k/x�<H�X�E���5�q��z��^2U�9��hfд�6��j�<�#�ز((�y�P��mN�۶�]����J�^��Wc��i\��ӱ(���?~I�o"��#�C�a� "���H�coM�ޟ՜ä/��p� Ky압�Aݩ�aO&��
�H9�3\*v;2��hv-4إ��M�3A�2:��m9�p�'�4	� �ì��[��R�Y}VM�oj�i�����R�z�R*��h%~�~?|"�|����)[�N�a~�	�����A3qr�{ž{e� Mfb��&4"?�H�Rt�%���?W6�]��ɱ�!X��~[���j�)Ρ^p(1΄.2��3S9Pjyg
^�KtY��šx��#�����B�)S}
9��-֭w�ޚ9K�#��QG�{���[w�&���6��Z(�V�!g�`����y���>���wV��*V�Yx,�B��G0VF`�p���HI����ɜ�I�&�m$���YAA��i�F,W4�jȎ�m�
�kȶyU{&�P�O(�DYT�����r���WId ������x@Yo�����*�k)9�_�U]��^�:�#�0HN8�����`�`�Xd���W�>:ğ��m���tH����<�^j=p�.GpQ�*ŶU���K��/&���q?������
��27��ߧ�l������LO����?�5��m��A�e��y�����!��Pn�/��3�	���<��D� �Or�I�d���K�p-�P��L8v���V�NO�������Y��	++�]�k��݀8�� �i�Li����FΓ�Y��tW���Y*�E��]�ar���F��R���,���S��<ů�v�1�y�M_&�	����A�xm��y_���ca�H&�묆J�G�u� P�2O�U��4R�|Ι;�<bL
�(�O U��i�l�l0l�ˌ�0���ASy�mE�0�T�s�ET�3���^���e�pXd��po: -[��D��F}O�:}�$�������7�~��2DA$��N��>��R'��Tl�/Z>���`���Q#L�am��N��P�x27J��g��m�3e�o����=����\ڐ��/�h��	Btյ@��y��B݌�;$'j*���d�n�Q*A�I��	8̇��M���΂I��M�Q3�}cG�Ƅ�Jʜ�.�9F�lg��C��k�s�w&_[ʥ�I�dh��ZK���`X^��"����q���duU�v���0dOvX:�A'��|���R���K��O������Ԟ����dl��`��VGg�cM��u�E��&�=a^�pPP�I�����I�[�qLѶ�G�>ȠyO�����Y�(����?Y9��Ŏ+��� ~Uo�v��x9�6�d䏈���� �W��茦8  �<'Yf�(*��H�^wꅇZ /SN�Yo�f����HhI�o��J�W�^��r��<���B��W3��W5)M��^d2�|se(�R	G8�p�t�����%C�Qٜ��$�⸢G�0��u�K�s4m.e�7#�f�D�f�6%��4ɠ��L�a�ם]\� 8겼3�P =pܕ����Z\4&���doET౴��-�R���Ai�Ut��Hz�-���{�M�Ǖ!ȭ�H1�.����>(����\u'���t
�f *qn.��	1!4.e׬��j�;�o�~;m��l�r�#�e�;�Ŗ}S/|2�R�4�r��'���y�� ��*ֈJ�Ϊ����C0���SB����E;��`�{,���I�fԻr�D��W�+[Gizɘ��г������:�]a���ǋ�<��[69��W=�[����$���W��5�@H�����,Z�]���-1S��]U/}�"dl����X�4�d��[R?k��g(�p�]�7��`��@�%�`������Zq�E6��� �VK�N��0hj�����U�j~�����à�K�?��L���#�� !=���~��鮦�ҙ�����2*8��u?�Vl-J��_p���Ҋ�]���7n��6@�{%��5��z��>��c$QVF��WlO$�ӥ6��ks��W���Y����9��n�	w��l
ĕ���z��&�?M�g4�um�Hkj�
����"�mf�3:7�(L�s�7$2j���O~��oK�a�e���w����P�!�e����"��`W�7�JL�pӭ�E)/3_5�/		Nr�)e]��V"g�9I�<+ɇ�{�U	��=��/i=|�5-?I�!mg���"�lR}��z
�[�\��L ~E��n6� ~��9�%�\B�7�T0G��K�yd�9�'�P�Kz��>"9^d��B=�@Zu����������'N�q��!]�g`)�`h�ǄY�'e��[&Hb��N�Ҙ��a�� �.���BG���ڋ��
J���wb��/���ŨEm��À���:�[��xx��a�g2�6�q��Tz �C4%�!?1Sz�p0=��X�����d��/G��t{z2D��b|L���M�21K���E)D7N��g�Zp�
Q���}1���O��7O����#c�E-嗊Xd��3�c����	����湯�$���1�I�C��*��Cd�[�\H;������wK)�U�3�UL�TV
�st=DLU/��6NdI�H��sE敼�M�%��@����giP���U�z�)a�Sx�P�C������s�=��C_������<�?=TJr	b��!�����J���;k�������%����\P'f�N=C�e��9�d�ED{��)�c>��������������>����%�:Ӹ*�벉7Y4j��2_�k޽�S_���u��A������<�kg� �ȣG��������M��M��&M����:yMU|�9�L	bIc��at��;�Vx�$����<�8�V&T�&�|��"\�JlwC�&%�����2�"��s;��n��J���,�8!�Cqî@���gk]�lg���\JIQy�$�=B�IŶ�a�B�z�6�s�����P,%t*�7Z��|��C�\���H��f�-�F�UP�3��o�素��X%��t�bؔVr��r9���`�+�А3��o,d�ꉰ�Iv�������>Y�� 0m��|��X�=�.E��lQ!�ت��7�I�2�;�>���͎�Q�H^kں|>n�n����NJ�H�����E5�\�*��Nc�Gmf��ݠ������Q��Ǣ���0�#��#~â^Õ�����Jj���E���f7|p[��XT�4����W�~���v�-�t�������8i{����⩳�����Vv����)�RL\�m�.`�sP7�����[WȲ��rt�9�sM)��Y���"�*�ך�h�7����C�hm��^�i�G�Sq��Q���ks���3��v]1������_����e5�N�뼩 �.1��?�/B��.4��q)�i�����s�u1Ea�<��3jߖ�`j �l�O�
��4׊p�b���0%�9�c�Yn4j���l��O����S��%p��5��|��q�,�?i�4���%{��d�\�S�����Ųρ�,������R�x�=����ƻ�vlauV��)��j�}�$�s\WP��ȧ�Q���ͬ0�VOrK�\]I�` ����)x��s[,v��n�F�t���)fu��ϟ���k�O�(S��n�����B0��r�iM�}5::~qYӶ���q��j���Xͻ�A�B)<K���,�Ppjdo�����| [������RÖ��Ә�*��v鷣�QHz���/LP�a����_�+i�w*����UM���RH�˧蝫;S�xq]���)�p3����LG�@�$� ��B0  ���?U�G����#����E��mr7,�k��vi����6r)�1��:l�1P�̱̱�fo(�g�e���r{Y��Rݻ2߅�Ksfفp�rw��!�e�<|��[~i�ͮ���4��v�:FlC12���<I3r?ⶑ��zW�Vвj�A��,���ww���<���ͪ���Z�(�����\K�%�`~��+L�0���jy���K���~-/�E;r��g4����+�' N1�$��ԥ���X��Z�ɒ`�>�	2�cb��N�z�L��D�]�`1�K�[�a�S�!�(�����$e��˸�=��w[R�a4�C�2 @-��eY��M�b���@�QR���P�ed�\Z�G5�U���]sQ��T1��DUM���Oqs� �,d�T/�Hk4�T-U����oJ���'R��e��-k���PlH|�sj�]idV:a����Q�8f��$1Ɩ��p��]I�w�Ef�*��-	�KE��m����R�[��8�����U�tt�GHǻ��u������)K�k ��Qg����%<��%���o�:V�&F��fs���\��v���!�C�p�W�Z�k�hO��M���S��B1��yѷ�t�͊�����ʛ�9��XfɊ�o*߱hnQ���V*�d�)��`I.����*��N0�A��/�7�2�*�l��_��7G5�i������d��5�N`q��z滠����l�ʕS�噘���r����K��}0�h���4��JH�E�>��z8�����'�&��5��ٌcE裮�g"l�4��N��("0�o���9q|��� IX
�J7Q����
.c�B`�aR���h�jp��Ro�{ֻ�v:���ΞbSfS�jwqYd�>��d㠿�~D�I�5�2�) s��܅�A���#z�E���0A�*����<����9��I�O��0��U���-�!�T}d��I%��Js��b�S�a�q#R����hH{�͍��+"���M�f�,�D�����ȩ}�>j�/�,�@d�~��Ӎ�?�ef\��]T9���ݒw�v*t_{s�%�Vx�����?M;��C���8�����6�X2���;W?���G�����U���L�{�#�[,�Vk͔�Wp����W�.ҝA�$Xub���pY,�#���P���?V�V#�!���o�g۝�"�n�Łں�K�qq��������#��X�� C^eW~2�����&�ޒ �5�Q�??�f��+JCYJ_V�~ؚћ�k�Yn��K�]�\`_L��}��.�bd	<b3k��Yv��`�
�<~�]'���u'�v#�]�a�<L ����{ֻ�k�U�,ŁQ�)��qa�|6*�0�H|��o7�x�r0���ѝ�3� �]D�L81 x#�"�ݫ�ƌk������2NM};��y<q^b��)G	�*1���2�$�\!k���h� �8��v���(���'(��雽o��%�ˠΉ{6��O�g�ʊ�o�u�HKa sV	y�P�E��2�|�C�D���PQ/�c1*R'���Ԋ6��i#K�����OG��c��6N��3�ҡ}|�[D؎~e:J�o�	��6jq�/�GL|r�ė�B5j��q;��PY���֨$���P�r�������ޓ��^�gd��zQ��ءu[.U�E�޿�+c�tk���:�Ѣ�j=�D�)o���&M�YH����j����0��4�սp�	9�I-r��r�6Y��¿�G�ݎ�M���z~�į�spf �y|3�\iW�U�,s!�N���I�
}t }#�N�o��>͂6��P� f^&���~[�	�4B����w����,�b�I!ߴ�x����}qto����������msg�����OK���^CO)�u̐^�u��&�`��3�����K��@�T�l��:�|�����I)P���M�>�M閧&�RY2hfIZ$��/4�����_ukA��-���2��<IX="7^��k��C��]�<�Ѷ���w��H�h�����f��n�K잦�I?1��z��ήu���Rs�M��ɃW���j��:Fπ,;^ ��j�3�~���Z�0n x���bqꍈTY���$oA@7=]�u�%�����5�F4p�	g��G"��0�]���J�t���=(T)!r��X���Vc�lk.�5���S<QLS�k�⸽'FG,%�ؘwz�����o�s�����Ec�7%�;�PEx�qr�����5�УK3��]��=܈5L�f�1j���b�g�����9���΄�%9B53��6�\�o0I9��"$���#݃^�PQU�47�uE���ݴXȶ���R�����*fL�Х6:�[(�n���@ ��2���Jb��m�k%k�՟]���ylR�WS	^�9�=!<��2�����we��H^�<]P���nJvP����9ݙnz�L�me����k��=;1���������kz>��C툶��ٙ<^s���.��N1sP�O�,�ԑ������9v@zSu�"G�}T�6����_8u�r򑆤y����X�
c�4���M�d���<�m5K�����o�R+�7���~)\�,�L��Ы26�V��&�ss"�6	쵝؈#�$!�'s3tln�h�@���&e�N��C�I��P�F�"��9:�%0�ڑ'gT�2���=�̲�.n�H6�C��'0��/�?(e���L�%�+c;)��-�eH�nL���'Ahq[5r�ԉob�u(�nV	L��d��M	o1����i���U���7.�����&0c>��=p.�R5$��2����9�)կs8�NcV8���*6��T�1k�c]��Yx��_Y�k�dQg/��,9.Ƽh��Y7ӚZ��\��t\=ǰ���b��?Y+o�/T�R�9���$ϓ�|�tb�P�m�.[�{М)Q��D�+�p|��z/�{�P�����aT���̬Gr��XY��1��,�0���`�Pߧk�����%J�A����jeGڳI��7�c�1�
������Z�L�s��7j���y.�9���B���E���wZb+�f̓@���
A���s��8C���ř��1f�J1���=-Aͩ�u����D�GJ.P�&;@$5:��o�*M��Y |�����w���	�VM�S�Iv�kD��ɀ�s��Iy���T����C��hj-�^
�eɜh�Tcy���'����H �C��jUj��)�&�S��3撊�M�d�8�J+�PR6����[r�ܕ��	�`M��/�hM��j��'Ӣ>&x���7lar��&9(�NK��j���~�>�\@�,q��q��Rʚ̩?5�߀/�š�UR�GOM�R) |aì�m>�t����$r��W�%��W��un���5��zq
`����p�Ve���l��Ox������6�A���M�[IԊsB ׍k�e��`$]a�늨���j��>�Dz�;�v����y��l�����6]Ʋ�7 WH�Kt�r�ur�7i�@ܩ��N�PyD��xo�c/a�L�֣<��]��_�.Z2AȄ�������Km`��$�(��Fp�M��8�o�a�!��v%��xu9��B)�C�"]��x�'Y�8���������ղ�A0�g�ZT��|Mg��x����������	�D�Z����ǝ�ۓwϵ�"�G�9�|�^y���nW�5����P�?�sx���H��ek��H�#	?���6'Pxӵ(���ɩ|u¤�z��Kȟ�$���e��������P��1< �LGW]b*xd����]�Y#��P����g�';^�/�4��/�z�x %L���'�
u�F-�£Dxz�ƪyaN~T\�+�5�g퓜=����+$�D��RU|����F.o�e��PJ�Y�b�_�쫋 � �9�c7fϱ�~�<�(����oh<ª�=)B��:B�j%��<��X]��$�j�	SտHC}%�d��q���W��=0�kx;`�0��1-�i? x��r�޽+��-��Oݓ�(�Hd ^���o�F���cB 0Vέ+N��V ��^4,�;�3\���=7��r�9ė���}���m#Z�J�(��gI\�K��LqT`�q���<uM�;s o�sU#����2_2�u3GUj;�rZ��͌���d�S�` �xE\=T��N�R������0c{����;Q�%��?�=בX^Nط�*��u��4�d�0����@	Q��sPN��J"�l>Փ�iH���%�f܉LI9�h�8�k���H����]��V�5� �\i���g�ݧ� "�ޏi��#"h]3/�8�&YJ�bwDo�,�a�Ą��K�@�!��Z:S�j��TY��z�<6�7��b�BbR&��( ZE��ҥ�6s�.s�@G�wڎ���Y�jZ�W����DHVMb�ko_��Ќ��W0���Zr1��0�#�[�N�q�0�|v=��A��׾|�-��]
�'��>�|CUn5�T���?!��qŪe3�v���t�mEjbi�`(|};����W�4#���j@�%�Ȋ��!f�sB��������M˩�Q.v�b��D�adI�E��j��{�cXҐ,�0~k���m@��7^�i�>��b�y���O�y�.�6DO�KO�$#*b6oI/�bg�ڽ�i�2f�e��2'|T���&k��6ZR��+��R����찰2��aw��e ���|տ�}�K5N6�"�7O�����=nG1�\�1�Ġ)���u?�|�.�o�/��N۰J�sr$#��rº@6��qǳ��Г�ԕ�s�n������>�4:���؜�4�X���׻HH�7��{ ɤkZ��%	)�C�K$��E��$�������^c�� z��#,��AR 	[^�['<y<�!��4��։M���"6�8J�'.xW��8~��O��q��4S���f(�Ө��L�-������h��U�n��	���s&�����S�-���I���r��̦��צ�$��n	��-��7��F���-�L�d��%%�t�_�S�;)�E^]C:�U0�>��}�g`���ԫ�İlt���j,K����2��f�v�4r���JB�D��mY9����ӛBn	&|�)p�Ce-5A�Qb�]����%�C�#��sV0ȥ	�0��7�<	j^ő^�*R���*��T��&Z�Eտ�����]f���K�o]_���舺��/髙��3��1����O�R��۹7^��EE�Ü1�c����5�.�Y4e�"�Jzp�"ᝊDN��#-)�u&���|e�Kr�D��+���e9�n:��B 2�&>Up&?t�;B�T�u0%e��3)�Ԧ�Ad�-����i��t<]S��\��r>��-HJ[9C���"��D�1�gJV^!�X��GoD�8�AP�ZZ�E���yy��hJa�?3�J�}�¦�pO��4�Ă[��梉�e��Iކ��#�/,�c�Ԟ~Ͷ�����{��`O�J�{%�!�R= �����B�̨-&8(
5?��Iw��9�	�t`�"x"\�P�Q�k@�UA���b5/�ˑjH���1||��&w���prJ���@�|ூ�K��^�x�l
	~�#�gQ{��0]��籴�{\�l�5?A]�['$}���������>)ȗ�!eL(�M����1��'�t���s�T�E�4�]\9�*��U�[�c[�*�P�Ac ��Uͭ���Ś'��@�d���F*�쬗p�R�p5��i��.a�@<��y$�q��F��k3�6��n��{	6.,5� �F;��ˆ:p޼���3j
�x��A��3y�	L���ּ̄6|}��oM_�͘��pꎃ:���F��OTc,��S&.�E���l�C!���I��gE*K�3X��+���5��x�c���B���#���dZgD�+�\�h���˗�k�(���v��f�����
���W���L�G�;C�FmD��*�N��J��]����GG���Њ�����:��@`�̶�pʩÅ����b�|N���0�c�|e�@�l���a_:�C����o{O@�U�]�����j�9j�ԓ�J6�E�6ak��#��T�����r�8�Gx+@��&=�foعeKaؖ#����I��lj:���`��F����ӧqM��;��&��_c2�"h�3��rMEy'�$U>�/vc����]E��k��)[���k�I��C�X2�ݘ��ʨ�m�[r��=hQW0��	��agؚG����m��{�>���9�B˗X���ZTnY����������W��*ʅ'�@�&�mn�;<�y�k�ޯ2t�[�I�Գ�6s� Ԧ���-��9�\�����_�0 Q�̨��4��+1����1bo��ϲ��	�ӻ7`�]S���{���=��A����#��\����,X9ǟ�<	28��TgZ���خ	u.�����	,T�m��>Eֱ*�ҳ�?U7�!�co��.�� '������Oo�|��GJ|	��o��8�C�U��G��;�O����r��[tBB�o)5����* a�^,���d$Tf~�t�4�Y �L�=~k+q�_�������G�K���-�p�!q�(#*��G#	晹�~�5Rgr�!d؄g�:��KX)~��&F޴���V�H���C��"@�,X�s�w�KX"����^W�b�r;4l��pݑZ�ļ��]�'"��Z��O=��z�U����N�l��jA%:MK9`w���b����Zb3�5��cey�%2A�:!k�6`��l�w�jżS���ˋ���:��6�S�gS�oG��#�;$���)�+�$Z#��2.�`�#����*�zD_���N�Z��Xd�x^�Y����Zɢ�$�d߯�*}}���n��VznJD'�ɲ/B����Y�	=R�#:��i�=:Z��_��JNQ��i�"�����0g��q�~%��OI'����]{���3�C�^��8�
,t�s�f�zYo��8�vi�ʮg]�d"Ƥ:�;�T��c�����E�AQ��}��:	�w���˪��ȿ�ky���e��\WB=Fv	3nW���f��n��M�ߡތ�O�t�6�t��-�e���4�?��x=p�)vd���tt����'���i��\@��n��e'sݘ3 '4��c@�!X�"��k�����ߪԦƳ��<�W��ge@�r;�rV�i�,#�n��h��s�XXV����N"�_���}]Ҽ���Ʃ�温�*�4iA0y���e�Jv5�kw�t���c4���H���.�!�?�j%�P{��`G�i<k6�����p�?z$(�Ãd���'��[k�{9�>2s���:����0�ʈ�&E�n|A \I{^�p���}L"�}�*��\s ֔�~�߿�v!�{�-�v�����K��Y�ϤO �k��e�<+CJ̫�[]�Ƚ�H������d���@*,�f�:�RO�J4��#y�������ɹ��<;�&3��%B��w����H��x6�v�r�;�Ow�@�J��`$}���Ǹ�� ��Y���#)f�踑7-��]n����x�,"3ZŬ��H���������.��:}ɇ`���T<8��5��ؾ�[g4�a����?P� p6a��G��Ny5�{�q���I�O���9e�8j���|�PS씹	b���CckޅV�|�3Y}�#pK��\���4� ��:M�cT��t�~I����o庋哋�e�B��r��"q'U��bK�-�*IB���P�a۱�-�py�?����S��*0%��y��t��X�y�N?�5Ή��\�`�O�jZoc��˰�FJs^�BÌ Ô�W�%h�P�,G�G�A�u:�	y��2iHb{���M'Z��q�qK�W~�-�pC��Q�(�U�(�[���|�)�D�)������R�n`1�	#iP��U&�;c{xɔ�b��Na�1��ޣ-�˶)^�Aث��e�As�ӓ�u>�O
8X0eA�)e#�����,����dQ�2o��͐���9�-����R�pv��/\�*{0��_�=b��(��f/\��__�kK�f�[/3T��!�ac�2�B��������q��ͦ�	r���G�o���x��sGF(^���eL�M�a�����7w}�2�����.EH�-3.�x��U���y�?�X9Zw�f�.R�ik���+Ӡ�AE����v�{DS��+�~O�gKY�f,Th�#�L���N��S�3��Π����H��2�l��SWg�s|��B4}q�Z)x�>�L��ɭ7t�a$�q8q���5�v�W`$��e�ɳ�$Á�Ru�	���$� ��
�o��H��3��kf��[yuPI�5��d�P4�F���F�4mRG�8��Q9�e�n��6ǩ��Ӿ4�\���N��ӪG��T���f�$�?<�
������ډ����3�F��$i�S�w0W�����^��$�)�{xlE�+�T
�9�c�{Ѯ8e4�X_��	@u���~t�̖v� wԝ�.��Ta��"|����3���s�'J��bI�M`Z	�_�_c���N���ή�-A���dJ�`w|*���<�� �=����C������o���-u��e�c֑C���]uo��wn���~elr�h��@���E�u/+�p�a�O� z��o#J� �T��E���l^�C���l����	][��4�q(R�hi��WqSK�$�e��F$�d^4��m���zF�r�1k[/�ᅢM�.C,~,0G�����l�lo=}Qn�Z�9����5\]̸dl"5km]Ee����^�x��hА2�7\~<���40�`��s�%�5O�2S��/8�l�u���S\�T��U�u:g����('�ι�c�N����dd���-�i���ƨ����c���&}�A҅���]�V$���q~�LyB��>���I�J���|<�k��4����'j������J���̇���p<��T�Q!��mw���7m�WF;����S��|[9��狏���~�qN��i^z5"b[a�d�v˩���w�<(��H%Y�5H���5�v���5�����Xz
�Ԧ�hf���&n��Ç�v2U�L*����F��Ś���,F�|�Ϗ۹o�0�$qG=y�-�"�MH
�1̆��u��/_i
��uo�`��H|��(���v�Þ�?������RN�A[OE/�p�vT�~f���v��԰�pu�l�O�/۞��Sh�\\n��=� l{0Ɋ:����$0��S4
���o������^��{ݽ�O����w|-��^�7RYCX�Q�Y�dz���P��L�1~�D!�	b�~wJ�'�\LaM%F|�|�(N<�G���Wb�+�j�a\�r�`~c;�9�����u#��t�ih�Z̊#�/}	�1n�����.�Ж�bE����R�*���j'�qr����-M`��6q\V���P�Uu�b�������u���`�2���́o�vv����f	����GcԠu\���4^@�������I^)r�w:��L�	��Л�YH[�!��s)���:�Z�Ǉ��]6}	fIB)�����n��[�
	���|�@cաi��K���}2,U��Stdm�����ו�ϋ�������朷C���\�<~�<�+��A5� *M`�������Z/T�*րR��Q�dH.L�5P�Se�F{��p�B���3���[v�LO�!P�T�Y�}������
��������U��U1&�*���Y�ƪrS����\��y ��9:�$oMr��e��y)%u3E�K�v�[[#���ηB�뮄��MoR+B���+���Js��
ߥ_+Y�.��r���,�=�W�hq�S��͇�i��2�M2���\�k�v��`~���H�o����hUpn?�Rn/�a�0`�7�TVG�q���?��}ɎW��� J5>�a�o��cQ[r����4�-~��J�}pL�F��08$�|j������6�(��%K�K�0�9��R��="NK��}����� us[�V1>�xX�ޕ'K6&�+t�5�:��̈́\[����nf<4���E?o�ͺ���E����d"�Ĝ]EM�D�>@��N�]~��E@T������c���f������+ğD���v!SN7�>4	�
���Ykt���cz��R;�Z�i]��{�7�r��$!r�f�M������r���w���|�{N
��&o�$Ls��^U)X��ya{�E	�+� �x�%@��+>������_���t��a��}Y�>���E���e���;����bw��ǚ{#�hV�_�X�r��?�� 9iQ�66���2�.��9>m�j��ǣq��K
'�<Hwҕ9�K��4~
��d����Q�#cs������_�N>f%��Y*E#�	\��k	�r���3�T7��vɥ��C����g�5�$� ��$�4j��=u.:�ui��M�����⵳��� Qf&g�m����Q��%�����.b�<�)���]0�<�	���$*�m��%8�����w;N��7��g��i�#�a�B�csoIf�d�����L�HLf'Vt�^�	����BY��p���M��G��	�!z��;2
���X��@å�|���u��K��h��V0Ԣ�!~�Zĺ��~�im�)��9�)�#lYѦ�r�\�T�T�r{�4�$R�e]�5ѯjӘ�]�%,�:�g������
n,g�,Y'��fz_U4�c<
���y��FJf	K%Z>I*�)W��c1�i�^�L���s�=W!>i|:%^�خɚu�NQe��SX�x�B��_�	�2Iв��F��p���}�v��6�J;��� ��S��Q�G�E<7Xx��
"�!Z����mn(��# ���y�gV�;�k�)q���5��|ˊ�ͅ�F�����[��t��)�P��8.
��l2�;Y� �Z�^9f�Ӄ���	:�R���%�����f	eG��-T����e�����J+��Vc]����C�ٽ���ҝX�j��} ����V�����\~��c9Vg_�{R7L���(�&'�,]B����of�a(���N��u5�u'��.��o���ml�I#�+<8����_XA[a��,t���|�p]�B	v��'�(>����ZG��WV甂����,������2Y\���w�d(/�*|�v��3��t?�t���`�.�Vą���I��!B�`���	��(�z;DnϷM��\��n3������$R�r���u��b)}G��U>�}�'�z,Z��j����s)�h6}~э3珕x�sAc��O�GWd���R��
�W���+ľ;� _GE*���A_��ϥ���͉���/�i ���Lx��N���9ʡ��B��xo���9�z .N*|Grt[GU����鈽�D$�WΟ��8_�� �'�����]Ǌ\�����A�ˉ!H��D�Q:a��M;����h�� �s{�q'�wTVy���s@D��ѐ��c����d�'^�Gu���J�S� �S�"���b�X �/B=/2��W���<taQxH0�8{u��C�&��šH ���(���lt]n ��5m9Կ�M���y~Ua���#gä���5�\E��H�V�C�j*{��\�ţ���F��3�o���̇:ϛ��A�}6(p��gY�h�����8�NB�-N�:��9�rqɗ(���I�D������z�@E�R�v��߭y���5������u��]*�'W�.K�Ϭ�q8,��q�Gw�>h�vsa�{�˰��
�Z@�)�(m�G���	�H�y��dʲ�\_��p�����_dV]���!j1�[FX�ٔ�b����4��e0��f���y���%ֺ���H�zZ+~��d�]q�=�M�r].�I"�mԫ(̙]!DH�_�a�]^FQ47�+��s�0�u��P�wbI02��ǔ�P$$i�E쫾�Ȱ��O���� ��֛�e%{Rl�Y9W{�d�L �Ք�v�6؈S���71�C$�]�㍔6߹
>����l����g�O�Ld�/�P�uU�s��5��D9�FW>=�������܀쥄e�$��s_t=�KU����𓋞�2I���.���o��\)��( ��Y��hV%L�(z��տ�?�����Z	*���C��wl>�1��rxE�P;}&�s�k\�5������3�&Y��&�}�i��cν@�#7+MXՔ>���V�+Ȅ,s[>��;���ax't����GG�hZ"}3�=l{�a�J�L�@�V��O	-0�Zq{XJ�W�nnG�P�}a,�{�N�"#zJL|XaL�8����6��+�"�(ZF�a)��n��|���q�~{J+w��5;ϯ�b����;��g� �#[�,>� [�����d�K��8�R�S��L��=V�(;�?I�YN�L���BU�]��pU_���Q��߳q���E5kz@&hEM���ᅣ:����f���lc��}�� �;Ek��rp��_ڌ>ևU�}V���LI(v�Vp'��zN���y�ʇqa�&�B�J��/�K ��VpNo�d%O7�YB��0b����{��oل�v����A� L��ϖV���xW,���;ux��6WL)�aC���b��M�fw�l����P�ALI��[rz�ku���+�����01��+@^��av�B�V��	��@�u�p�|�ֶ�I�%�f`+#T���*�c4�hf��;-Lb�/B#&���I���Ŕ!.>���LٕWu[�u+�[��dOC~��4q��\>�N~��3���lE��w{W)|�]u�mӜS����f�M�$�>���"4�KU�8k��}I�(K�����㷋��uB����SaZE���5m����2�u����/��Q��iY@D�js���`$\g@k�ʅ �߈L㘝R���X��,&�� P5��·X�*:�f���U&�7+����܈�7���N�w �NG�3`©<dO$���@�(�Ħ�YW��p�U��lH�����-7
���jq�:���������L�{���9�By_BD��5H�\�G7��+��w6A���6����a�W4]c�uU�%k6�N��M�4iZ���OT�:/��4�exބ�X�&-��2~��;��K�1��l" ��S;�� P�j�S�/1BJ�T3A:�a��*H������L�~n-������1�E�nl��r�nb�b�}�[<rC_�z+�E�Al�N��v�O60��9q�%X�n�l���(-�H��.J_��������T?�Qa�=�ܯ7��`W�'�0KS��/�	yj֥�L��]���8��[�_m�� V�V��ӈ��]��$�����e��r{R�Tt\ǃ�v>@���Z�]i:�7mè��nɑ�>s_��҄�r�i�F	D�Bqٛ1SU 15pg����_â�-�І}J��>X�	�[(���
�E�:f��J$R��w*����Z�RYT�7Mg9��)��������m��6�����6�����U#��54����]cΨ ^�{����I��fn� T�g���PJ��.~NSgp5�w�xhZF�l�� �\��r��v�U��´Y�& �����'��F�[Ӣ�\{AmG�l�Nv�O�{{{��$���d�8u���\4>��z���3�����C;�(�Nt���:I�2����Z��I�J����
��<8��":�.���l �fO~�k3�n>2Bt��)����[��ڕ�Xϳ��Bi~�KD���#��<����J�~=?C�C(,u;)�1���n�U�������V(r|b�ҝ7
Eu]��vBLŮ�y���X0�`�^K��$E��J�= �5�ˤ���1Xp+���]L��*%bk�}3������%"u�t�Z�`b�����T�A]s�dcL��u�l��q^T��
�'ŗ^�L�}����Zh�Vˣ0m�=*���>k�#2۩�1Q��t�Nw���	��^zmz:�Hy��Ȱ/3Mfc��2���SP@bT�����G4 ��4)�o�a�s"�k���y|S�D�oxM���{+����ݮB'������2�}X�0�]�S��D��cd�[��t��v���=�q�{h@g�F?C���Ʃ�Tg�>P��>��@09�a��{Kt��Oյa�����#�Mo��"Qc;ލ� ��3Q��k?��A����Q�����%��C�+�z�v���D)�iC�H�Khc�C"�ˈ0!�	� o��
����6��t#x�\h�}z?� �+���	N�z�q�?�eAjE��f6�L$,�2�~��ʏ�~����`1I��h���o� I�Lp��f�n.�u����R�`�Y("�c��z|���D�1���F�'�Y�?g����	��,�;��X!��+����^0Q����(Im�OS� -���Q���x�D�کʊ
d�Y*��ЭL�3@y�>W+��'%������L8 �Mf:�z^�U�%0�%���Y�viB�v�ao��yF��UƝ�o_�&��� �t���:��lj1y��7��&��@Xp�Qg��Na������
�)ץҩ]<��z��K�x�k�u�YD�JE�֞���x�b�-�;�b�jӘ�щ�B�&�gw�S�
�3P���%����=	��3�Bvo�\.eE�'�B����M>�6���V_%�icQ�a�-�H�؂�g���Db겼[��4/��E,��e1���-�ol� <��>��{B�땫S�b$�薲�%�<!�"��X}ԄJ�����(����H�����>J.&���h|�hc��dø�~[Z#F�u�g��f_!yO��+�[04�04aᗾP}&rM�� � 
�I!v%$q��YO.�/W�P�j-"�+��|��BD���M�X[�,:d�4�9YtG�2�^5:Ō���(���o��[�<��1KЫ�\�8ڰ?��C$���EeK]s]�VQ�r�?�����[�(���R,����"V;<ↇ�Td��&��H�A��#�AD��Im�+��-�20_�>`yz#��hw��|[m1���g\1�ԡ��)N'��R��Y:�*ʲ8�,�I�w
�W�eԽɠZ�p�4l��Ua;�_�����̧�Bu����.�'8��x��P���}���Ú0Zy8�1|���Fכ{ƻ8@ѝ6  z��"��d������|��#��d��f��p/V^,��At;���(IT�������X�dh��z�o���C�g7�8�WB��z
ai=���M�mcԋ������1~J�!|Y�w.�F��ZδLyK�	|�'�T�\��M��w�rS9q����ȹd�>���(���aVg)�]���`�#en>Qښ`�!��e���x�l�}�]�V~JE����?�	β��Y.h����S�b#(.��i%Qp�2x)���x.��$�B	ʚ�8�ԧAx�8��m�#�u�u��s��]��
�(����c�?^w'�9��P�T�r�Dxc�g3�w����A�9����F��b�p����}^>�K�� �\��>����|.��gc��U`�I $D��w�|~����!�(�ߨ��j0{�d5;O��H�#๸0f�^�Y7�!�m\\f���"�hm�8�,��N|�yB����y�4,"��uf�r�):���
'C��g�Vn��^h����l2����G�����n����>�`�"Yi9R�5�CwX%�U�j��#O����z+L��B�f��Z^���B�7�T�zLA
�L��n*D���s�I2P�}E2�5~���`���#� ��P'�#t��Z�����Ȋ(��@��M�H� �d�uWQ%��b��m7NG&�-��`/´?�U���\��Vx�+͈Vdx���e+t]��lЉڢDk<�����.U��1&��"%�b��%��yhVB	�bJ���C-AD(��ԕ���م�ӳ``Y�E9����p���~�)��뼜Ztj�Ef�o[�H����,�]�����{�o>S����/��~B�>p~T7>C�Z�~iS����&��J �֯��,޻�]�}x��2K<qD����살�/����OIB2b,�$F�Y�{��"���y{��\�x��bYypS��7��>w�����>z��u���b�pq�#"}2��Ta堷������@s�'�#g�j�C&���@_e�Q�y�߱L�..��L4�&�j�YiA�وe���KO�Aa�'�@����4��6�S�I%rq�۾�^�����Q�X<���9+��F������:9�S�+�ȡs�X��Ҟ�?��Z���~������_�X7����^��Ca"�?H%�eY�<�HJ�OfM�ZF�W� ��͑E\��}���'���-��7�(?6i~fwj)�u�ƀJg*vRNn_�b�􌑑/n&�ى���3�=���1U����Ō� e�P˄�H�b���;S�<�b����7��@0��PL|(ZX�=K�S��?���l)p�9��ӑ���o�߉��j��u���G���f�t��́4.��K�D�#N��0�ڃ�u�heO�uO#NR�ZO�R�f���q�e�4��3k����f�Q)�_6/�F�U�t���)��q{�h!��+�eaS?z�����qk�R�/L�Lڋ"�6!�c�w˻E�03̼��Mk�}�����B}�v��\,+>�;�ζ����_]��Ʒ�����f���WM!_��a���9Ȝ{0����t�nYY��l-�C���}z�f�����:�P��h�����t>3�.D�/	E��_){�#:�d�u�:0����Y�1`\XY����ǚ[�]�7����n%0\���o���Gz��jV˴�,N�3���rd��e�D����CI�3$��Ýa��g�=~�q���Է�\��s�
���5�E��
D����L2z�fQ-ή��JL� �>V;�+�H���(&�C��>ǋ���� ��=�h��~;�H|�^������,i��&b��T�E��,&A��>�9�T��V�F&Kq�䄭26��(ɩ����9<���7l#�ou�M�+5o�n��{j�`���=#�n�G'(�[�����,^Y��V$����e���DњE�x�;��.�h���U�;�N�	q�Y�c��I�A��v����k�ݵkse/=��x�*�B�j���ً������c��@~������* �>�=���c����m����Kb�X���M�S�'="�7PD?��,���V`ap ���~�7��y�·�Ub��m�|dPR
�Fi�	Ζg�:���|�G�Y��K�(|��!FC�����᷃���G,iv�=��L��(i���6.�Em�1wX$1r����[n���m�uȶ ,�5��)�vʸ�3���uR��ho�x�_�M2O3�\�IY��-� ��v[�k�D�3��5�IBm��M�>f-!�7�|y�Z�zϨX|�'!G�u�ק&���f�G���#I
���a�!�)$7�6o`����n����3�l�j	�D��_6q/�ڎ�@������J��.A��V�p݆���f�d�A���3��'�{�"a07�x,Vy�yw�MA`�HZٿ7� Ca��!/�~�֛$��-��ky�}�\�V� �2�}{�ǌ�n�ԑ��	�]!*UBLp[�\�t����B�m�S.���{Y?䛹�X�,`R�'jƚ�f�V�QV���n֣�ֵ���\� ����z��+ѻnZ�I�ӕ�o�bP����`~Ck����Y�0�� �>���/L����0<���|���{)�ˡ�ټV���;,��sG����[�X�{��j��[��ߥ�ԍ��!rr��ۈ�Hv<���`bF_~C�v� �qWaب���N	�\��7	Q������h�*R�b�r����]���k���MY�~���+������N,���6����G����n.%ￚ�8,p�r\��:�5����S��O1��m�a�n���;���r$�^�	��T�|Wp坾
H���_�R��E�����CX�G���n�j�RK��2�'��q�'�|����-�����J���;������ ���4/ʖ�喥����O��]s����Ĩ�^ַC��PO/��k�v�H_��Ԙ5���T�u5lh1�=%�}�r�oiU
1�eOE`����U~X�l�t1D?����oup5\��j�6Y]�.���txh���0�v���:�
N̬��>��cWj���8"�{�j�(є>*f�@��C����ϋ��̩�q7Y��jQi���(׊�5����zu��Ԍ�5ș
�<��'9��4I�Y�P2������:��&�[��~Ė��SXu���HqM�
fj>������2P�A������~���3mt 8�E:>�B���95�m�N�����R_���Al"�p��e �j��(�zS�@p��"��	���ir=�o:T7�{�D����
�C�h.��!�B�hQҸ����e������,&��N�w������}1Ȗ��
��_�Z�ж�����g9��|�^�j�P���?�)[��)�:���N�q<�����d�;��$Rs�q�%T���'�C��;z�#��f��w��e 2j�H���$׵��ԇ���6�b5A\��3���&7����҂��Z�e~�(��%z�,�ڬY��%@�m����O��.�T��T�����uD?��g� �8��Gi�P�C'Va2��ց!T4��Q����<�����9��D�E�����|��T6���r� CÃ;���Z�[NǂkU|�;�oуɏ|Oof֎�s�TI������z��7��55F8!�q�\㩰іc�����1]f㛋V`4�[:/�tLW0�f�a
K]v^�F#��ettR�<~��ϢUyR��@�e��@UT\�jcq������u9����:x(���VT����vR�v�M�`L5;�(;�9˦�����V�ţH�ݔjq�[����S�%�R�����IƭC4S��ޤ���1�6�x3�< �H.NJ?�.~!��" DM��u��d
h����Z���\ȸQ*?���i�K�s��h_��.��x��)w
����b����ح��[YeW�4dٹ���M��D��,U7�'����6������{���K�,e�2jl�S҇���{Ӛ/� ��+�$��]a�֖Gc`4��W ���moӉ�|�N�b�ܥ8ݑ��n�o-���=�L���.��m��jp{��Y��^�]vz���׭V�;�ד�/��$�4�!`��L�"7�Ŏ��`�^ӮY�D6�,%?X&��Eh+UL(��Z���ܹ6���F��B��Vhk˸s�g��N�*5ԃ����@�B��x0,W{�x���Lq�Y:�
Ӆ�s�@�<�X%���cQ��-'o�9�fE�UNq5"��h���P�{�P�^��P�b�	��"�l�@�H�����{azI8ށ�΁Z-�S2n�0�š�s��������T�w��b)�|s���x�_u�l��MF� �W�s�L�Tm5�g�����/��8=�v���� 7$��W�A>o��+>�� Uh����@F=�S/7���6��3�iضS�`]r�N���P��J+�:m�Ͷz�p.^�LK\�Z�,�*r�N�e?��\x�
��h�W%+�-�{�������������b����:}l�\P{~"E�rA&F�� 9�c^���C5��~�m���'��,�b;��C�y�?��2����� Q��v�;��
�&:���w�P��Ě�m��Q_�	�\0Ô�m޽�F��g�Нo��S��6�u���ѼƖ@����<�����V�Р=w3�֚Z,�M�R���/��^(0f'o��m���YFki�g��y�~�����Y���m<x�*����<ٱ������/K=�p3DA�>��]�p���=��� t�c��T`�@0�k����:�+[ɱ�����b�47����b�9����n՟u��dWp��Q�n��!;�'�N�6Y%SWG��Cj�v��>��yk�E}�l�0�wrn��A
;.�O而�ot=�P�ܳf�]@���@9�'�!."x"
������$7������z#�iՓ ��t|kb�2@:��Nhɘ��d�f�X���7[�с�gxߑ�7}��}N���{Sb�CJA���  ��w�,���IC�Si�Ⱥ�C�;����%�o4"فA�� �t�r�T��D��GNHf�S��iD��Zi<�S�GuT����3�n�y�և��]��f���UzA7{�vT=������\q�IC��i��߳IiD;~�]sbpX{��� �9��oQd�\���BD̨l����&��0t�����	��y��h�j�H}1����2W���a���#E�88k�k�8.!�L�؂Ul��8�L���n]
�8z	�`CA�����˼����� �ȩі���$�ͩ��`Ɗ�c�J�4P}-Ah����j1��Y�51f2J���8;��ۭ�&�O0Á�q,��"L�ϩ#���AОV�����q�L���ϙ��t�@o�b��;��������3\EL������~�wa��c�.Z����j^�ʝ�\V�����̯,�3a�I0wuH>�����c���s��N�`KS��k���&�)f��v$����ab�A�;�[T�w͎��~c��[��<-ƻK~<UL��&��=<�TjӞM/Y9����Vm�Y������i���s�W�l����HaqH'�aΣ�weǆl�%H9��F⼧ͭV�>� B���׷G;V,�)�R|�b��;j���T	��}�%����䜅��v��)����2��n��RG��g!���P*bP����F�=����U`u�g����{H��{7�[YP����9q͘k�P��>vO��H�޳�\΄�sz	!�e@���%�:�p�������0=�=#r�4}�s�D-ݽ�	��[�&��Y�fk}uҡ��P�m�nR�P+��,YZ�^മ+�4t ����d�D���hm�@�{Lʨ��]4�τ��h.���zQ�w��9u �,�s%�6_cH���P�I��Sx�-F�]q������P�!�I�=�8u�� y��X7�0��H߁ϊ��_��O�uG\�0~� /W>�&���������g��y��dp��(��0�8�pPc?�b�ɯ�a~�2U�ҿ�"�gAPS��Cg
�=,Zc���S���f۰V�Н���K�p�������u"uQ>؇��J𘈶��֒k�kkX^�ބ*�RL50xv�� r�@6LTe���IK��dʝ�- #-�C�>�sq�,@�����Wvi阀!{]���Rk�(0�j�O�!���u-�-�yZ�K�*A�yo(m3�4�FRR�ps��H�35������:�c V#" ���c������f�нY�!?6b��+�-_�}=~!S$��Lz�T�ɉ$��^l3u[jk�ܫ�
����j4�	��I>�n�
ӽ�*��w�{N�K�GT���o!^����o��z3����M��c9C�/Ɓ
��E�?�S����0����b�jn���&+@�bz'u�-���P��+rj�Od��7����W��cD��_��J�~MHOQ[�^b�]�H���D�H�����5�5���̖Q�����B 9�>�y�'�.B����Wk�F$��rK�S�C��)x��l�
�֫��j�y>RF_�������:��T��PbM��`Ԛ�{�L_˒�<�4q��D�D�aDn��9�$�>P�����n�D"��g؃?`�4s�!8l<��cq읈�L�	��h��(R��%/P��?I����E]��дU���F�:���_\�`3ǜ�aW}1�a�,������-�Y�=��̹/E)S�u ��O��<H�Z�bف\�nJL�}
p�k�Qj�*l 
������A�DLb�u*-���CJL��+��	��ZP��f��:�2Z�`p���0���L��cmQ�L�΁���Gi����S  �aH9 #�p���{�s�y�� �� ��pu��ݢ>��ff�����T�w�}̼I��X�	�����%�84���6�Am����3��:�ҳ\�8>�fy�&��2���1�ݚ��.UC,e��xC�V�*��D�O"WjV��Y�c_��6l^1e	��
ք���,�0��.�����d7�ZХ:���~�a�\g���e$�]�z����WT�WH���6h��֒Z���Ϣv͙�a��xK����TI���e�����+R�^h`L��𿜪U��1l?�d�����6T0*(��U�N2Y3�%����9�Q,�ع4m�({��������-��.\Z���%�2N���k�wG������ ,E���^PFrS&C/&j�q�b�i��m6��ZW�Ua!0�=틨�~![��Tenxd���yʒͬ��4e��0�K�w�$)�L�bȲ(���!��$�ɤbιkZi)�L�R<�\�O�X8�9���NO�R�U]�lh��ŕ��퀾h���
'[��{"�Uy}�>Ax��- G�Y�g��Ճ�����9Tf�Z��d��� � ����9'� ~�a��4"�1��k1��T8� �L{�9',cM����f��=�j���!_[	��|�R�_TO�o�Ĵ�51���h���HHc��������.Aphn$Il�R�*-������,�X|��qŧ&���<M��>_m�c�i������m(U�*I�;ʫ�����@����*�g�����������]�&	�
��������q���b�|�;����_�M�
��|7�?�F$��&���jr�Ն�d|o�j��_�B+b�ങ��ߒ���"���\�B����g�\���D�:X��Y��ز�jQ�sv����c�����P׵UZ�OT�	�~�|x�"�$먇��;�>9V����k�m$��F�����$��o�t�	������(\5=^D(��B��$l
ݿ��n�4�*&�7ѝ~Z��TN���.�ց��J7�+��=���I�q+]����˕rfE2q��}�s�w������fp�x\�'�#���e����ҏ�$̓ΰ���SO�{�G���Q����h��UW�G��5�A\��o�L��oZ�����������J<�r�tq"��d�h޽T��n
�tO��Hic���b��pa�i���vD���O\�� ҍ�[�z���~�rg�����WȪN�8���� �5��pL`�V�Z$V�L������.��k5���%_5���{7SPt�.܎�pxQ����n�N[�N��Q�S?������u�-	7�~K������"�Ǭ��{+̵]O#��|�:/RS^�����k.�7v��W�9�Jo2�h����Տ�Gό�n������Q.X���vB[s�����_�U@�����(��Ȝ�����n�y�,.���6���sa��J������IG4^�fj�Edo���v0��P+|=o&vP�X�!گ9���@��L7��#�T�.w]BQ\%�Jg{����-���2�G���4�~���]�M�j;��!L8���	Ϻ����\]�gs��`\�z~V�Őx�{R�˂�B}D)��:{�7� �܋��d��R�5W��^{.A�ǎM�@'#����=XΦ�j��{�m�^ϴ��Ⱦ'*ߏ���	]�!����PE�	�!n:�Do���WZ�),�8��L����YLg�}�1YA�w�4������A�|y�[�nwz�;��,η��K��c���J���Ip����+�'l�@h~@���N4u}j�xYu��P՚뒙#��'�Ҩq�^`���KS�3i���ҫ��q�I���㌰v
/pz��!�T5��$�a��]m�Eboz��G�rJ��LIb^�f�[�x��l#C��v`���X�S�rN=a��
>��/�s<�DeL�Bo#����&h�i��������Ca�Yh�Z�/6Z�F�#9}!���a�/־���8R���I�>�ʴ{��K����}��Uy�i���ւ��d���Ԃ���C;s?�8��r@������p�a��W'���	����������lzꒃ���e�}'`)ť���+�bt6����Wn%�ҧ�h�ÅN�n@�wm�=5'!�����3+N�IY� Ti�#���iY��|���趢ͭ#5��\�U��8�]����a��胦�q=�U��>�Qkud#����  x��DX@Q�G5���¹�CA�rE��y�%�$@�VN�����#W����P�2 q��Ы�~����o�2�[ A�<�X��M�����*�٥K�l��(��B�ߕ/&�V�����4B�?,�RU���������	�x�QAoO��Բ��+L0��s���W^�1v���ͥ��940'|�nGqQ�w�2��3)+K�\�5�GNȕ��(�Ѻ�<1�8l�y`�O�qM߶'��<b^���5)
�wj�����U	�j<?{�����}��_	�-G`c���&��L	*���&� ��F;�=F��v*d|�iG)�-�J�=Bi�����gHO��4�C�`y9��k��q&!Y�0��NŞZxh��jj!ݿ�"�K�2�}���I�i-��3�0�#��}�3�?��V���i��c��$D!�4��W���C��t~��i�a�����z\	�(�+�c�7�5��[P��È t���	0Hu�^�zY���J��H/VR��Ic��;���@�Uw4Yg��(/�T]y`Α���=��V�6���t�ÇǖE��v���J7��P7J̓ǍE�������B�X/���j/���&}����+@���2�w�05�/�sQ�'~���8� ���J�r���vA�[���S��:+�'���u�'tSǲ���H.��>NM"X̨-�_{���`E&i J�܋1.���Hw�-��٤/!��-��A.� ��LS5Z���˂8�,>�Q�����a��o)4��fz�=/�m�ܑ��.������ +�V�x{[��(��n>�sw���8�O=�T�;����p}Yyؖ�w&�T��%����z!e�eRs���	A�8�֩w��VEsÅ������N.��@q&��ۃ���nR�V���S��y� j2Y�MU��lC�y�Ϣ*�q�eѥ�b^��T���{���k�G�rO
�w�@&�U�-��p�A���U�$i%�vO
 �e�vDTT��֩t��6�y6�!%���>�>��U��ٳWom���)	��Z���*<{H$��:�>Ph���E���i�bH:K�q�n���ͱ�CI�S��D�$�&�ܺEdK��WB#3
�{����EqEi���W�=*�ޯ�K;�a�e�N|:ڿ�d�^٩I���h�`� ��lX�5��$�d>�ɸ8��G?�DQ�FF�^��f��HĶ�����u�Wc��� ���[r��~5)�U�j$5Q	�d�x�vw�B)�LҌڼw-��(�����qAc�0��&��.[T���<�b����X�[$�.3��7�x�ʨ�S/�Ӎ�F�ޘ=�>(��P7�?�DAhW�I	Xy���$d�i��ix�aA�c�a��������qGg��
$v� 3�l1���~�L�s6'�ާ1,.������+�`C����|���j���~���o=�u��}.&햦eߘ��򝹵��๘l�PFd>*�����u\{&�F����,$qrW�?@�m��h~�������<#T��b���NF����tG�1B���Vy6\�(H׃*E�:����gC�k8�Yj�M�A�a�S�/l[�FP�ӀkT-I>�9�&�a�I\� X�`c�Ć͐�l�l�1� ��^1Ŗ��\���^X��e@���O��O�Fp�v��\'Lr�I�ˠl#_� S��R#t�f�>=u�Z���3K2cf���.�����__W�E<+RHz�ɷ�X3�
�"��.n  �
~���DP����)���txst* I�X���I[K�^H�����a7�zF�᯿����%[��4�4��q�Z|O_�Nե�T[)�^�g�C�,�?{\��ŝ�\��>�D�ies�]� ��R�+s�j>���`���������r�>�Wp6�o�[�WD!OLG�N�b�mOGoLc��]�n�o���"���i'��ic��d'�#>NB��P0#$�,�.嚤z��7(d�ؔ܅�a���m�L��d� ���<='���!*W�=�Z���8/�C��j�@�(8G��אq>$Qe;�m�}5�#5 �>3�������*p���:�nZ��%�c���3b�]d�mW�Y�n{j{u�I�������?��q6d]�H��{Ą��a�@�}�o���-�n���@���v֪�=����1��2��c<�C����ts+)%$��/L+^�ai,�c�Ö~��M�z/�2�O�>�c��	!����989�Vo{��dB���n=�V��S7D���֩������`�[g����=JQ����|[��9]���/kkQ"�]DO`�P�C{	����6��O�W�NI�h�H�������>�(�(�*�C�8#JU�} �z��K|����oF��%��;rZ���h P�|A�p�+ЧiBaj�t��"�\��v��ˎ�~��_���f��\B�)yV=<��1m�
�l��{e���}���c��t:����+������Y�E�� Y"�䰩��]3��Țp��(�OK/.'Q`�I�y��s�<��ת�������o����3_�x�d��`��|%��Zp�`���E�Ih�!P2�A����L�(���"f�a�+�&��6��w�b�p	����?������"�)�nh������d��dηOњfx.j5iQ�k�+i4eB0!ڶL�R�k�Nk�dO�^�9lߜ{��ߚ�ot�[l&���Λ ��c�o'ӇtE�c �)�x�|O�U�X�O�l�.0��w�naT�k���������!jS}�񵡒[�t������������}ώ�i"bq�N	S�u�Yô2�n��Ĭw3��OZoJ�⠺��7.t`GE��;q"�"wv
��Ǜ��NC���p[Se�$�T��m��0�n3���w�8�:��G³�'G�,
�4�Gر,���N\����;Ҏ���]��:r���u�Jji���� [�����|d�cV�b�����О4հѻΤN���zs0����V�T��`��?�>�i2ɤ��N{Ĭ#XF1����2s�RP����ckP��X���\ں;(��Y�I��ec0�}�/�8=#6Ve��`e���m�r;�V��3\X8:"��ZV��]z���/�/��%7�;ԧ��U����P�t��|\ȫ��0����ӧ��s�鷪9�S'�)qKh;j.LY�xY ���F�&���L3�-���Z1Igy��n�:F�ˆ�k�϶ܮ�����x��+N�ݥ,�5x��(" #�1Po��1,:��5��)yO�};�~��v�j��ӆj�x��:{I"i":T�`	!����d��6P�t79�Ede�mK^Im�N�����[>$��f�ޜ;�{��+'O�:b���w�۸�n�lƅH�MV��7DH"d��7e�,g�ԗ�]}������=H�/�'J��4n�E�2s�ƪǮB�`�64e�hB�\O�����y���]W:��-\�te84��yR>�7[R�s�q�!]������+�J���6���|�o吏�����w�q���<�m9.�*����~��ֽ>���,���z:����s"�ׅk>�T.��4���ߢc�ql����EY��,k��o��l�jck��P�H;
]�����*�7Q�8B���hk!�d�W��8��BWv�H���L��u���6Z*Tq���72��,߆������
e3zg+ �\JS�C"Nx�/4��K
N X��V����Lh����+��uv���5 ��Qf7i��"�f4u:ߡ@�/5ڶg̾	���^*���2�O�]l�Ą��`��z�/�Ι�^����3�B�������Cȝ?��_zŝi��6ix�x�[1_L.�P���j���#v+JoK\�sJqG���}ΆG�l �e�^0�U
�E��˞$,l�zO;~�#+�;Ǧ��|2�*��w9�F^�7���u�ה�?2�E( �CM�#錑T��{j�K?o���Yڰ8����6É�Ql�j�tV�d?4�J�H����T�a������z؃���/���.az��g��~��ߪ�9V=��m$K�^r�כ��e���1:x:��k|��JT#�H�#�6b���H�M��u�x�qjR臭�_@�^�)	LdY)%��m�Y�� �y��=s~�u����}�W��[�W�������φ1�n�o�p����>��������`&e�8e�P�m��"�uU�6�@L�4����[: NT"����\�Q�_Pf/����䀫֨��o�8pT��Şܪ|_w���aFޠH���~��@�Օ�`yI��o���?����E.������3��V�L+V�����4lqm.+� �k�)�;�$��~����5r���Y��~����ѭ�k��QݨIf��8I�xP�o�th��X��a���o5J��"�>�q8G�XڱF�N��{�+�<����r�1�K�C��I��;������)����#=Y��{��L<!Ǹ5��i֏�}�;�����|:�uKS��g�f�c�c7C�Έ��.j���im���v�� S��}�-�PN��
�D�� ��~c��{�z�H��M��D@p�"������iU�$�8�>S��5���y�h|1 kn6�DG��ݸ���p>
�wr����Z��Z}GY��U�|&���N?f.'Y�q�ѻ�T����$���l"��ռW����T��0�Ԛ�H���ՀR$)8�ٔ% �N�OA�7�Nl���t��I$$���#������^�m�}�aYf+�c��2�,���>�8e!���*���@�˻�V�;��@���;q��	��0A��G�o�q:`�>`j�p"O-H�w��5*G���
� ~�|�w� �L��}��-��,�F�gt�dV�]��Ig�|]��ݺ�yR�K�N2����{~��_^���J����_�J�߷����(\X�����q�r2^a̘�X\�lb4���VS��Dٙ�Z�DsV���PN"�A\��������D�/I�����D�~K�����|X�dV+�����e�itR��!1FRD���λu?Iڙ� D���6y��5�������q���+zJ�@��ӝ�2�'����긬C�X�l�z�
���qo����8���8Aa�7DE)�Y�O!�#��,�^!yR�� 8n�� 3��txk���4'�o@9����W_����i�(��й�N{��'$��
2{%�H�w�!�z�;��gp�3m����\ňx��L�>m''���ǣ�ü���6���6��,`mU{=%��H��T�pZS�� ����zf�(��8��F�T��<1$v_͕�0���ڸ�z��7��(y���� �����̑̋��,��f����#=Vzr_�ٓ�;[�!d��}�G�߷Ę�m��n	s@���UϦ
�4�
	ّ"B�zPNK b�<QQ�yn���R<���xG�R��}o��^�\Ё�����ۗ*���'���U �f=$l)�]�w  ��o)�r��T���f�]0����ۉ�e�e�7'$�W�����1=��>�A��zP�?3#U$�B�����z�z�B?���	#�|��+���B`a��Cm�/����V�{I��F���F�Fj��RU�=������xߟ����)0ƞ���|A>��Uf�;#Oے&q3��7� �|Cӓ���x+&`z��zyW&L���?����wY�s���5Y&���+��'�Sg���լ�W�|G�J�)�6`8=F����G���mE����d�wb���W:VΑE�70�d<o+6au��``���֗ ��җp�Fs7���͟ʉ-�[%G�Y��f�G���p��p���1�s]�H��� �i ��S-5y+���"NR���׶I��.��K"��sY��0�>ŔN��1$n;rR���5*�b2*����>!�kݫj�p��)����5�c..|���GG��'�Q߉T�'P@jl�׻��5��w�c%t&�"��J�@�lnc����y7cf�J�uNURk1���-}�Uqi�����-,�d��ߘ--�Ƭ�zP����,���㨄���M�N��|X�գ>S�QV�ޢM��$MxY�-�n&cz!�!�W�I�(�d�,��U�lx�p�` ����)�1~W6	46��q�!���Me!I,��b��-Ѧ75�>�r?yl��
�W�Rq����*�E���G��To��:'�3L�vk$RB5D�Iz���i"+J�`�M�t��p�t�P����UVߪ`�V�W�`��@t�5UBV�Z�Gk�P��9��u:�{�F�C���].�i�'C��c��dv+����j���u���f�Vٿf׵{Ĳ�<������YmoP�����V���s0v+l��`��tCY��ͧUːC�	sT���.��09;�!�����[�|�<��7o1k�JU����qn� 4�Ӥ�]}~'s1�����ܾB��V��e�X[�5�6�Q듄?6����h�-,�X���j��PҮ tsmz9��J6�6� je2��v���N��eY]���t�����(&�Z��ٝ�c�C}O>(�CL���s}lDC4t���V���U�㷜���t�D��kX�����#��Zǹc���D���m\�˶[r{a�٨�C�P#-A�Y8j[&�9$�
��:�zB����}E��8 I}�%��R���)2� ��F��f΢���K+Fk<���&u�~~��o"��F2���i�� 6i���wU�#S������Yk��-���� <f������_���W_�O(�3Ƚ��km�<�8$����[>��k�T6�=�F��������87eY\����"!�S���r��H��.��9�}�����w��A�(5
�؀m�-�򡦆A:j��q��Uȯo����@��G��|���*	�Q5�qL@�K�@Sp2�����9l�Ƀ�z���������
����L{�0�9�3�Z(�|��Em�4�Bq��᪟N�K����#	��w���M��fl����R6SW����e�=����v���+�����2w�1o��9��P�nt�y�f����A�m���A���D��0��|.[3�����v�?����b�.�X�<{�C긫w�#����ݐP ��F�*^�[�����)��r@`���`�W`���ymIe9L�2g.4@���>������BsX�Mz�g�����>~u���T���c�[�����|�C� ���0n:�/WPW!rd)D�<���M ���Z�'Rα,� ����)��C�����*�rc���HΗ70_���w��S!�cQ�K}�K׈h�U�Ӄ��rn�� ���CR{�SC�N�/�p��x0�2u�y��)���͟�}Hk�Kp�+��s�@ l����Tu�F&��)�����Ĭ���GҦLК��p�J1��@��b!=&9j�2���gC&�7Ȟ��x
x��i�\;�xn��ʾ�Y�,;Tּ�Ug�Z0�`���ӟp��'!�`xi�����q�>���p\�H�:I��GN�d A��g}�J�U��٦��@p���	zP8(���{�~��ON����cfE�T��9�SM��:�FW���|��}�F�v៥S#J�_?X/�㙶�s+`��˯��!�Ж��|&�^� ~h�5r��[2�%�9��j�e{��"���u�[�Q&�ʓ�^�+y�2N����S�V����5ݥ��~��D�dlG7�1f=�>-k���\��k9�_b.�P������C/'�a!�O����u귥�}Q�١��<�xP�]�c�Z�V�Z�O�>J�����Z!�nJ�T�n<�쬐��;'��p;F����u�:���h�ͩ)@+�//(�2�"TQ�G솙�4ZU��ܭ��]�����Q���_zԴHg	}F�L��Q��.8J��>�g�l�m��-��f����WN�m��"�N�;�Yv9�tC��:��[�p6٫U��r	_�kMO�2/���Ǳ�_Ԡ�"�V��e6�],��+ŉ�u�`>h���	�����vEd}l i֏�NrM,dp����.k%7 ��]����{�~8���M�z��x��$&X)j�_R=���A}0v��Dk�0�������S1���p�?�9���bR5?I��nk#q�ݞ+޹'$?��])A'&H�@���ap$<�,�>tm\G6�-2ۣ�f��w�m�Vs0���5�K7�3�;��{I��G��C�k�����"�c�ႆ��_��>G��LK$C�7�r|��� �ؤ���*��u��x��CT4��X��h��4�t}�ۗ���ٍ�o9'���\����O� �Nn#� D�ѭH�!�X� `���؈�=/ME=��������s��H�X��$�(��h�2�]�|@*��d9!<,��w�r�Z���JH��\d#�[��#� Ex�V#��'2灷ßnB3�F�*�;T?/�2xpI<rV�"_ϷH�"��NN���gs�3m#6hT�J/^�k�~�N� &~5��qa��}rO�Ou;]�y�b�W����%5�7��DVGh@v�L��v+�.4#�hѯ���j���IѢ�v)P��[s���g�����[1�7i��<���v]��MOE��f���\��	�W�F�
i8n�����Z������Hh:�+�����n��Y���Dpұ�Y���*'5y���;���n���E+��]��RiӒ>o?h�y���mieT=�f�=�m��7(ޭw>+��� �pNd�,��6H&	1=Y5(d���gB��Z� ����y�2n��u*H����.������Ȃ�ؽ�l`��IJ�"}�-z�/`�g�P�v��	��ԩ��b�T�t?��ZUa�Q�a!G_='���M��"ni6\�|5�(�D��l�Vzx�?�`�"���0֙v��r�Բ�PO�x�]f3	�r�Ig>O͇��������Qn�����.�5%�jΊp�!a=�Mj�{�W AZ��M߰�C�Q��)Fw��N���{�?�vA�P�3KFE}8�Pކ�W?�����k��T�Q\��)Å���`3����/�R�Q�0�~R7Ulek�?���Sb~��	�����E�d6����h���T� �tэ�Zo2��=��栠�����/P�y�.c�������}gVw�y����M�~QR��r�6!W��#��]�6?�i4p��ʤK�X�O�{�H4z�M�♉d��T�M/1�J�q�0�D�> �EDW_^�-J�Ƞϰ`�yY�Ńj�^�q���<�Z�����P�9?#�,� �w�\a�r����u��טJ��:��y�
C��G0��~�e[�����N��(�&ذ��X���y�3��R�C8{a�J�p	+�'����C_9�y��B�zb�* dl~V�Aϟ��?/��/�f�@ ڻ�8����6�c�n`��ݹ8E�6M�d��$� ��S$j�����,�IGvh7��?�fpm7н�3Wu�psq�7	n{�2��rm�j�N�x��^�&�}{���n�����cA�����ɒ����V>�4�	/�߉:V�����o�22���1fB����ᗌ��$�^^E�v�I{d!�X���Ӫ�*�|iR��j���	|.�&D�~'�]΋%
@��0c���}����3�Կ֢�=r�q�s�@m���5�|���[ʃ����==U�v����ݻm�BxH*����%�x�����P"G�۬�'<��0�]CM�2��R�*y�?��7M��E�z"��$E�����;!��"Ɔ�]�t��x�5ͪnU�s�A����ףŃ��&	�]ѣO��`D�	��8oG�U����ᰐ���t���uUYô��Zt�"���񋎆�1�����O�D��ϭ�E~3�����[X�~ܧ�s-}&� 0�n�`�v��Y��CU4�&�v�2V)Q�����o��I�\�(��y^+���/y�֥�_-|�Rm���'th��91X�|�����.��_01��D����jU�ʩ�A�]���BE��B`	j������Q�č^yB����o���-��4�Fr�2w.�F��Y��W�x�{'���Q��f�_0����p3P&��e�qJq�G{g)pi�*0��ܥ�'N]�)��7�m1U�c]<P��ߨ@��ۚ�&��!�-� *I%<l�y��P��)�Wa�X��T����:^{��Rn4�B���3wO�ғ����ғ�~76-�&��� ����_�Y��/�줇�Y�DX)���`���h��*�h���T�����N���(�����Y4�5��>s:,��A����Nj[T���l^# �53��렜������!l*ZjIGW�U�N��*Jԟ��8N��ㇰ�aLJҀ,]�<l"<K��zW�G;N�$�ነ������)(:!�F��F`Ҳ�:�G.�)B���E{�Żdl�X�2R�Stz����
F:��>�o�\\ޛ$�{�ws��P�E��ODn��q�Wz�"fH���Ў��8�<�5_k��U]�p��8���[N+O���f�W�2�]�o�&�����7�og�� ���+����/�L��?�7����hq
��rf��_A��Ć�����1U`�_��o��|46�e�_�Qx���$1���⋵���I�R7� �/�����7�������S��F�S]�^�%�ͼ�A�(����m�96%`�,$B j�e/pc��Hu�77ú��n���M� .{�XF]�E����D���Q^�=/S��\[UD���J�05	��==�����:�P�����)�]Z��E.��4��θ��4�n2&~\�wkF�\���}���ub.�Zw�����$�f���T�\ZTNs�%A�F�S����f��y?��8��xo����`��2�gw��DPrT�����Bx;���*���ř�׬���;�Y*�[��3�k��� D��>�:��]�t���
��=�eg�[��y~?��h:#����|O����6�aG~��x�{�����*�T p^�pB�<6�urC�������ؑ�g2���S'|aʷ�(N�/6ZE,v.��zy��a!�R��Ou�tREyܒ�D�&M��{^W���X(���}5��|F|piȢ����u�s>�M��q�y����%r��E�-D}����Ǘ�Ď!p�Ɔ�`�qGv̐��jb|6 ��!s�M'5 �9ME��ȸ�Gb�'q��p�a��x�Gp,TR��]��x�� |�bn`F��9���j��Zڳ�T&=p��5Z�)��`�.9@u��73�P��_^��߻lӶ����}�)	���D���ze���إ'���T���
4j2<b�p�i8�b��!�O��Q�`�f�WQ���'��6v���IsfJx����<���'��lt��RrR�Q��b#1Z��β��er�צ�H��.��{{L�U]�XVb?Q�i�vq�#'\l��B,�5��;�s���y�n�9��ӣn���R����UD��������)����t�hH����2ݡ�|�A@gP����+!E�y�>�g�kЖ!+=!^�O��[2�eR�Z����Ic��r����	#e����Lo�0<Sɇ�1��ܳ9�M���_!\�ZDo���3�"����Sy/���@r
	Gjr��V��ܑ�C�j�'�Kq�"�9<X� @PrVw��yu����H`\o�D���h٤N�~��AU��7��s��o�E_�c��y���K�ޱ��q��۱��[B#5�����ao���G���	�j�H&�Ԑ�(����@���-'�z�ɂ�	�r��+��2���s�t�LZ�1ƶz��&����o␰��b�{ϗ1� E�&�ew��e��̃(>\��z/�:yS;YZ�	��" d#s��^�Q�c���81�0�BR��ϸk�'�F4Tk�zg"t�u�/�˵�A���1����q¥0�/GB[�!|������b�+]��T�3 �Ph��h�޹ �g7����{i�s��f�#
pq���e W��Gصϑ��,,h7Ox����W�\R�N�I	>R���Ԁ/���tpo\9��Ϳ18sB�.�#e�VV�x�T'��k��oH���¨�R��w��|��/h>�hb
 �K:�ې�a�91J�i����#�3c��?��:K�ʗ������{׉:�G�� ������Tc+䩡�8P�z����������~\2�Ͱg�6K5p��h�_��,�%�p�j:f���D����-# ��d����!rvj/���?�N�W+Jq9��i@��F '�F���lD�?^oYЧXIh҈���r}2��2��I~�z����[;��/���z��A$댒#֟�m�1��ٶ��_(���_��օVS�����kL;	�ʔ�#�E.�w��J6z��t�[��J�NX�k�i@�H���Nή,��a��{����9����J�K_��Ml����򕫔��w	z�~�l8D�G|�'������_Dl,�|�>}�b�����]\��!�?۞��Skw7�:q���E��qjbӁ���鶪Fn���n;H@1�jD"45�G�YѼ��b�N��?*w��[�	���QѬ���u9��ؐ��Ћ�>��!b6۞�8�z��m���иDKZ#3H0X��k�;�F����N��:�Wma�"K��V��:A]���R�����<�>K����%q�7��e�}�f+CDH�=ƯēG(�M�iB@La���ZQ���l	��5}z|��M�j>�l@%���A��氈􅒞�iԭ�5�2({��˽�*��\��Y(����W�Qf�>a3%{pk���%�*YV��dg�}7�<�x0�&�`�@EԨ��.=|x �c�8�L�V�ȂVC�g��vة}��4%����(M3�/1��g��@���5�0�����Ï=������z���^��	澑��aDE�<�����9���49R�;���3i��
�#��
���✶։_N�׳��k3 �Ӫ˿e��P=�W������aA��;G8}�/�4Ʌ[��i��|4��&+�� +^|�����n��nX�0��	=.b[�No�9�KYt`����
�Sk�&���4gQC�������r@b�ȗ���"���vR���S-�:(������(������v���A��S쉭uH1�	\ 9��&��%-{�e�M��%��i�}4B^0��=g)��̞��|_p�
>�=�[�5/�%��F[�~��&)����OgӸ#�%.z������;���E0�����0�s���,���|��Vv��y�5�Vz(~��`�� ��hU\�)�AΖK� �n!���f��������a���0���m�;.ڰ��t3QB}����ʹ&=V�'1���^�&�*J f�.�k���uo�YnN�orpR'Q�+@{p���6�"Jø����m�w��h�j��g
�
�#q~��ϔP���9nhrS��LB<�_�|˯a�P�hx���/n�kY쁝ǽ��U�D׷9e4;�7���L�MX�i�l��'#j��9]�����`뜷�wࢅ�ِ@�.$]-����:�P;�h�
��@��	YZ�m��l�3'b�-*z�i�j��.\��8�
�����e=>���=xā$���t2��<F�T�����	�-P%��͍�V:8>�dp�JB�E�����4�)q��C�u��S9<������_�ӟ����j�M+��N�y �PHB�I��P�E#)�8r�;���\�p&*Y�4����\�l�o%�Ҙt$95#��Gc2���3/㎒~��Ucc������(��]y���oȞ�tn�䲯���?)�������kD6��<T�J�K3�����W,j�����L�6M��<�y��2�x����o [��5�h�&�7:`ą��]��4�VRE.�קt��N�֦^�DE;���@y��X��c�m�6�2W,�[�4�%7�
	��Y]e�������x�8!a�kP�gad�=����6�\�f��j̜8y�y2�QB~�g��r{�ce$�����Y �BN�lJ!�
vJ���v�#Bf�OƢ���Ŋ��_58%j�s�	mj��M���!M�_:��x	�Q��IA���J������!Հ]���D�Ў$��7���4�<V\�#[�">�×ys4)7�u̿~�j�k{�������Op�l�'��fI�O�!
)��{1�Gj"L����mU�8�it���_�U�^L�<o��L_#E�6">GC������܅8�y���I:��{M�/f���]�stg��-051����A V���Kr����6�̢I��l7%�eR�s�J����-�k��)�!Z���6��b�/?�s
�y\Gm��c6O�'����� ��-Y�)L�Uq�d��0�������"�����E��q�g]�A�\ `y���9)U��xT�0�mt�,q�M�!R%��k�a�M� �{u��R���BV1�AJ�ƌ�2�i���b��V�'�<��T����[��`e^�f��D�G�G���߰%�D�1`0����h�wcjM!1i�{VN�N��ͻ��q�>�`�7œ�ANTeZ#y�h/�d7)�}��}9�~X%v�� �u]��k~@���V�L��?����Z��s5㔷�����c�N��׷e��n{�B�o��<b��l"�!�Kj����(nfr� �����9�9�Y��RW��e^��a�y`�E���,l)޹}Y��&?���^����B�E�(I�`��$$s�+h�J�y졛Η
��*CJ_1n32Ǩ	t�F�y�廀���
���\�ˡ=��f!�9�p����>1�fE�X�����k�#���o=$�����w�yy� ;rp<2(�F�	ts^5�]���_��J�2,���m�� �pI���֠#���0|��T��V���׸z��&���%O���p
..���Μ�䳽�����\밳����գ��:��1�_���vۘB��G�|9z��Ӗ�ˇ>�~�f�y�_�9��
K��啅ok�����޳Eds��	�A�ЁgS��+>������Y��~�CF��}�n�S��sJӦ�zy�ut��w��.6"��龄�Ɣ/����#h�� (�Tǅ�@�����0N�(��n2���Y��Y�H��N)��\"�AejH�|ݩQ�tnA�[d�8�i�Gr�7�I���W�y��O�N��jW�����S�>��:��fA�����{��'��n�a�!�f�iN��AL�$ч����^sL�tEg�5ސ��C�����"�C|�yL��}|�_-��?��W괌E��Ż��h���P�2��ܮ�NWN�S3x/gsZ���6>\��hr^���M�ɼ����$ʵ{y7 h��"����pLwt�t��(yʧ��s�Y�k�<5���`���[����Î(rÍ2���|0etVk	�ҫ�ɤ������&-�@Q�2�w����"x�͹N���1���O6��ϻ�8~>�H r;�=HY���F�~��ϝj��N,�R˛�)��&���>Ȟh@�c����/��I��)�@�� 2���c�vM����R���s���cl��ߠ*1=��c��ˈ1��'X�Jf�~��Cq�~���<�������ΆX�U�Ĩ�8�E��]��C�9R�¯y�g��◠����p���UW�H���hu�'(����G���\�u��N_�0�����|�Ӵ�"0��6�.G��]�ڀQB�fW֬�L��m�gN�%Cy�7�>Z�i����PшoܠPW�	�}g�OW�_&;˚n�miB+���Yz�����N܀�����t>�� �ݐ
���j���Ԉ�k�<\�l���:�T{�M�蓍,��Dن��Y&���N��}5���0 ���O���!�مYbf;���&:!nS���� K��Y2F���z��<�Jܞ�ɡ���fV��ZL����.�	�Z&����w�r
q_� #dA��7�=y�X�ϯwk�Qi�\ȫ�<�w+k�*M�h��ҝ������� u�lX1��c��Ʋ@:�M���5k�ϨB���ت���M�E��Z�-�Ԝھ��$V7*5s&�M��h0m����b�}�72@�q-6��^R�c�\6��+��#qh9��Qx�)�]�7<���c2���p8�|9L���H��?I�g]�܉�q�R�ً�`ˌZ1K��X��ljm5Rr��ˮ�; 4���u4���X�J}|�cJ<���e�t���IHH��.����L��`ن�L���(��<wk�W�^��@����*�'֝��Ǻ4��wT�Ήv���퓶]��� b��U:�9oZ��N�`�.��8�����gq���j�s�ݘ�շ��[_��s"j�>ֵ1����[�Sy,�6[t�uFi<&⾋�4���qG�Gu��Π�E�e`��ـ]D�o��|��e1�7����F#��nF&OF��ߢ�h��������ۘ�2����O���n�&�f��L��~g�xt�W)ό(8�1��C8�k����Y�H�+�^�Y�R*35�#`?��2����SO>Bh���x�<A������>Y��B��� ��"0�A{)���X��&xH�i7xcc7	�8�y���[O��tc������jRV�0R��k� �#N�^h�3X~�v���)�aLQ��Ν��Ew#j�0LQ�;O����E[9-r��F�������(����{���'D� Xni�^�6h�u�Ee��BWŐ_ �Z� �X̔����+l�2�IXj��A�vv>��_�w#��ߴ�{T+K�����e��/ȸu���,v� ~b����s,pj�b��ϛ�g����{�Q/��5ze�F�
��P����3m��mmxB��.�iZK6h)��������'���ڔ�7�R�A=7+gw��U��������uk�x7�a��&�!^/*{�^#�P�wwH\�ˀ[��#����Z�r���L��l6{x�_���=��N��;ʕ��U�4sՍ��ƫ�/��a�C�Q���á����������QA���1�R��X�I���Zp;�� y�Г�Y����H�~�6�&����`��8�c�0��}��y�	�.d�8~�W�R�~:� +ASg�]%����x򍒄~�,�,��/����+>��X�5��{� �n�]�G�����M%���GRXǵq�Y���������br��m��gF' �L-�aŵ�d$�V��|�EC.�6G��{��1[]��������$�:# ����<}%��y��^`��]�=Oz����)�*t������j�E�
�����Q�X�o?��D�����ȍj1�]�`ImXU���)T��1��<Sj#��,�$����Z�CذvƠ	J$��%i��F�UYP��44 ��Fs�>7��p�T#%m?f��(C4$����|
3��G?G3]%Պ�W�������ʽ0���4ȵ
��ԧ�ƶ@�S��G�����%P�c��H������,R\7p��o�|��<�3�����= N^M[�EUc��K������Qy�Wݻ.$�l�� n��V],���@�5YD��C k�X����"���
�ǀT��G�������`~��~N�cj���,�ï��L'�yȚ��,�>�HlH@��d�vIךvw$��Ћ.������pF�;�5������U1���QW~*���,�dvk��U}��F����@�9*h��ty%͓����k�������@ ��ZZ�8���$>IHtO��e���_�v lj���Ң�]s�#�e��7G��7ݩM�>��=G"��?��yT0@�%��]��]�][�T5���M�k�hE�z�7
x���8�ѝ���mU;��Hon�iοfp��x{5�wE�y�m��N��-]ttW��<���g/v4��v<2�2z�5�C�A@�]3y��g��{:���բ ��A_�o�r �m���e�%�*"�����F�An�u��<�l!'��,�P�U�Mc�'O�1Їn�`����O$�i9s��s�b�ڰ/�����l�`����D��p䔩7�|n!{�<����N�'_rlC�h���4�ϥ�~:�2r�U�[��t����/׫>�S��c�u,�}�B��r� ��s#�v��ѽ���f��ߍ���r	�Rf��'����
UD_���k���򬛁� �ǣ{��?�v�n�]3j�����#J�Ѧ�����dD��C;:C�#FǱ�wC5� -�k�W�0ȡGk0������K�<"�7b�^�R�9����|�Z�(�qF�d�Ε~�>#��������>�6Э1&�p����"+����R�fe�<��f���r��(�Ӑ�,��5NĨ��<'3q��|0��8����"2��'ARs�����\�!�ޔ��"�2q�i-!�f6*�alM��79�N'Jֳě�P �j�F2�m�*�%�x �*�T|T!��ޗo��,/Ǣo	��#Ӧ�_�U��_�]Y�:��J|[m�S�������i�ȣ�V�)�}�, ?�V���/�FR���-��)x���Y��(|��V詖)�bV��"�o��jUOҒ	pΡ�����1�e�<6^�ft�*��a��w� p�Ӑ��.�"�]zgF]6�:�LF��B��N�� kS=s��	gR��늰�.6N�1t7]��$̣p�7�ly��pf�q��I<��·�;5TK�w�����V��JC}z��&X��D�$U4�Sc�">�)�u"~��NuYk��9��J�%��X��zs9y��K$����
:��粭^�u��H� 
�{��SUS�/@��rX�D��,⏤E0�u��7{�A��;3��*@�nY���D�� SM��O�E��6\�
�g)�������%ža�47�i<r���円�e|�@t��9���-��O:�/gN�7�Eo�Eb�vu'h�k'*��8�Zsw�o{~���`
{2qc��n��~�s��q��<!�����/X�OJ�K;x��a�NE<��z�����J�ݿc��3�Ma=����׊j�gl�vt(�{w2�N�La���@uqpMHs�}+��U	�������� (7��҂eS;��� B�j��
*!�T��.���ë�^B�� z$OU��\� A�`��܏G�
Oh�	)Tn�6��Z��ѳ`���x��C"��5v<]���e�o�"�ܹz�c��W�L.�Jҙ�(M��U�9�y#M\%{s�eŬ����}(i���a���a��?@A�d�kE�z�{g���
� �GrU�qI��c���V�KI�@�t��B���2�|�-���o�m�� :I�:�9�ޒ/�܇�^y��7�A*�Au�do�o��M4?�>>6�qvA��������%�Iu��l�ۓS9�P�[������j�TAN;���pJr �Ht��bR�>���1��vxN8�Ep��\�߈T˛xl����uN/�\96�4`��v��|�A�=rcj�h��!h�bbn�IbK]�`{U�a>�� �&��hh�I� �3�Iͻꌑ��O��k�w`j(�[�v���m�Gi	+��3D|}��r&���"�]~��"�lr�3�zP����ǘyG�ӷ�݇��3���?���|���XUת��\����꿚
Ȼkf��k��������ʑJ��q�|��c	#�48����!�xZy�#ƻB�A'�88(�-�4�wp{�>��Ս�HA����mm|�-��#��6�DD��2���:��2Dv,����P�#lDS����a8�K�*�➜_!i�P��]����h;1v�1jSÞA���ѳ�p��|#-v/��F-�&�g@H޻��T�q�;j�
1��^e�]��o��/�H�!�4xI���ൠ*�W<�av���s�q�%��_��vH�_0&cF��D
K,�}M�
��:���x�.���Nz�RE�U~K(<b|j�X��v�v�ps������ VW�H�u��o�|߮�P2텆#H?����v�(n
y�&��/� .�Ԋ�y~*��̈́Ԭ�+�Yտ?ݒC�sn�7a��ta��":�f�Y[�R���q���0�z��v6a>�%�ͤ��-�j7Ȳ�~-4��������$�0Ы���2�H���%V�8�X
T��BMg�u�xB�U��X)��ɫx��@���$�)o��R�XT�r&�����&A����t^%z1}���G���a�ѓm�#&23ZqcЈ�h��y�����������)N���B��۳0�z���&�9@��K����*c��c]F��B<%}n���\ڇz��gR�	ۄ�W��p�����W�����v�0��w���C���|x��1O�F%����خ��g����<�mT3�O�`׺���`��Gi���Y��������1NZ�N�%���6h rQb��nf��S��rCT��z�a�6W��J�[��B��[L�mk��?��j| ��7�w�=���1��![��C�N����l�%wD��a-DLafe��u���:%R��l���Xv���X�ږ2���5�L[$�٣[�+�AJ�@��}�=3��z���6u~�*PS����0ڍl���iQ}-��2��g3#ر��g�gp3��'ή�O'2�|��/�@�ikr�
�q�W���)�G�o�RNg*^_�fG*��3^�}"�ۺ�:���Wk%����\dx����+|<�y��*���Y3�\S��j���-�5v7��R ��z=��oH�z��%���F�t7!����	��cGL���~a�_L0��и�L	�h���� aִ�&�`5���(�$
��]���aiz:u���g5i/�}���w��[�v��#�*��#�N躁2�SU�ڳ�ʏ� g؎a��Z<�V[\-j�u/���I\�~^ce�z�(�!�y�����V$s�6�DZu��[�ȕNXtm_��b���~�HO���	<6ٻ1HV*��,�#��y_�������kr~����|Q��N��tao�/�U:�[�_�`0��wD��]�����{o���(��3���~(FN_��@�׃-v7�����|���|/c[�XF>���� �|t(�m���.<}�� \3s��F���()Jjщ��i�Kl��-��R�b���5,^�a�$f��ܱ^<�,����e9=q=�v�^�SJQ�2m�;��Tr�<Ο��,�QK:��6.P����1s[6	r�fŝ�t߄q��x	�D�nU
�AH���DjP#`$�?�ߛjY�U{1���9���N�^kld�徐�a���8Q�k��À2�!=!���tn!��%<C����_�Ű���	o§в�7!�]�8e�ܙ�h��j�?���D���o�U�Cryς`S7Mt�G""� ��Цh��m���g����ޣ`�R�/���[�E����|�\l;�y�ʑ)��a&��1���J��9���|���L�cR��E�'�j��a��'q�����k����	���26��5��Fl�Q3�����D��(�9~�pb�@������@��q+�>FErRT?~OeQ��<|�ȅ�Jl�V�qZ�M� ���+�W��&���<�����~���L������¶�]C�o$�d��R�T��-�𪠯$�#�kgV[�a��r{-���l]��c�� �~X0Z̛������
��T�������l����
�B���4���|@���%�ً��T�]���(����I�)��
�>���{Gj_/}߿�TL����<�������/U�|��bK�?���f�#�����Fb�^M�64���6��x.z�l�1F��^ޚ�*+H#����
�#�aBg�x\E\�L���o��j����);E&�c�p�8�e&!���7���� �/�l_�]i1��� %8�b�?��<]1+6�0�ⲟ���J�%�A�r�(H���!���0���َ\�x�����x}��"z	�P��$O�e��%Dδ�_R���j�AV�\���s��!����,�8>�;I�k��R�8�ۇ1(�	���>2EU����@;�T��sUna�� ~sKn��3����2�n$�%т%����h^�2���)���SP����[�9�iş[~}�w���!�<�9��Y�>u�A �T�əVSV�c��l�I��C:/[�s�w��' ��|�%�W����=�q3(2���_2��x4jo%$�b�rVmf�2P8a6u�O�;��6\����k�nQ�w�2O$���(����4?O?0��Pk.��Wp���1�2/���[���%^���!U����tS���'�bԔf������CW��\F(���;-=����oG����pa���#�6�f�l�H��h���u4J����IZ ��\,��8`�-��Ũ��������L�y-(bd�z�]�_[��WHR*l"=�F~Emz#'|M�r����i��8�h��
�/�d-:`���)��O��i���>ԡE��L��}�$�Z�����3:]��OǸE����|�'�p�GD�	 ���Rit���5E!���i���OW_��N����F�%v�X(@|&\T��T��,�y�O�3M{��Ro��ێDn�Jb=�@=O�㼣,��+ה3��G��J:y�o�ٚy��O�X~�o㆓�FiW	e4Qs�J%�"-��^���8�a/k����QܐB�Z|��N��m�*��r��#be<�����Yu]j����(�k�W;3�����R㣻�����4)��D�� �z��V�҇8qv�&.e12����z��.W,��@V�D�NF.��/��V�`�h��sߵ$g�$������9��閟���9���M��NGC�� ��ZxR�&��(wIjf�ݷ�&S�C����m4�>��������1�n�H��c���|O� �o�~�r�=�m�U���!� @��"b�|�T}x�Cu�8��/�Hb��\4�����'����qa�~{���w^Z�̵�@��w��U������e�0�:��K���n"n(B�v>&9��}�����{�u����X/D����2x�|,څ��'�@��>��h+d���}�ٶ��5يA�����Lvjp�!�e��d�P�,��Cv��^�b�
r5;Y@pã�z�!����9��E��.�;������.�a�<��N�^H@�$�Im�$�{�u��#�6�(�N��ִ6����T'I˭�fɱ4}�/���"	
<�ː.]J��!�.�uX��v8 �4�3f�K�Yi6Ţ��Ȗ��:Ǒ����L�M�\z2V�i�J�;:��Z�loQ����d���MoB���S���5����"~UHP_/��t�&h 
����S-m)��LlW���c��Rn�@��.���0�T��o�F����hF�R�2(I�N�Ǳ:���y�ۑ���~^3es�iL~�D_N�2��o�N�8�5���<�=޶��VPSPo����J�6�y�N�*jC�����r �|\�5��ZϗH���d�Z�~�:�H��M�f��GMc��p�A=ZD�F0hdr>.( ��x�	�NZd�#L�E���S��=��b�v�+������6�;�ȵ�O��?X���ܼ�gx���-���` ����Z%���"��^��XC�=���xfR�b,oK!2��M �$���-Y5�̭�$�<b�m��C��2�����\�O>�m���A�t���B/�륂>��D�~�1(���ߑD��J���Ͻl�8�)��P\��,��p����Iͪ��}Nؚk�9+)�6�Fu�׎|z(I�NvK"4�n,�� }��d:�R&k�����6jueSJ*�B�Edt6���:$��u7T�R-yqL�|�з�V��Z�G���aa�-��������utd0��ͨ`�-���y�%F����lg��ҥ�g�n���s!��S��o�>p:V`�혉�����yZ5��u�#g>� �0֣sT�)O�t�m�l�
ϧ��\�Z�aPQN֡��ӱX1$�S�A&n�d*)�r�Acw���~�� &%��$�h�*Jb��5 ���G�n�Gr��^��X��J��Q�0�3�/Q��)O(��a�o�(���%oU�����/�t��m��A�k��7�6��Ek5����p�t]���P����)�3X�p$��	8r�G�XqwAފ�N��Z�+K��ޗ�K��b���1ĶBd��v�R���X5�%�� hd�χ:��j��޶��)�q�: �}$"���K�X6� '#�,�yP�z�W��Xq����#/���CҢ���k�I�'x8��gE�r�!�o:RmM*�ƋJ������W���	j]�zvI�#���u�N�m>�����B���(��L5B*S���ϴ��
��A���8*�yWo���zE�u%6 �Kq���u��8�Tc�s�|����������0QUr��`��������,�ǩF�%]ϭ��[�E�li����]k�&s�������a��-D�+�2:�s^�������"s�;���VS������W��b���������Ċd<�0@el��{&D�Q�8�����ͅ3T���kP�y������,����zg��C`�A9�O�������}Z�^�,�"�ĵ�o�!�s�:Vk兀���ӕK�ެ_-�)�W03��z��]��b�j���4�xl��S��-ί�W�4/@'����u�^� �T���-v&����0�D���}ABٳ�e�+H��Ac�v��(�a_)f�t�:��	.���~4����'�0���Z�F��,�4ӕY�K�9���>M�ө��Q^C6��wW�8Z4�xMr�X���βIi��׀
dvE��ﰫ���K��j�̿,��q헮�E�Z�D����/<ݐ�.�y"MGz��lL�f��jIo*5��7����Sq�*���N+����Eq)Cg���>��@�*͕o~�[e�X��P�,}�cif��?��U!��x�L[^e�^��O��V��1�쬶��W�e}mT�_-�!��P���j���Y�Iz{��b>{��	�_�ʫ��J;�s�u���*���"�$�C׎ڠT�`�AE!��+o
�b?^Ө���E}!S?�O�BR2�T�6�N\"2L�8�Y1y	ݴn%�TV�`<�߈P����|%@N`_q�	���Q�aT�'Eo��rZ�_g�9�ӆ�6jW�Q�0	<Zʛ�e�o����d�V�ZW�7���S�+9"Mqd �����@���2�s���c�=�W����EQ�֠����z�+D�,�\�����K^�~چ?�nf�fv��BC�h
��9�f�I��
ǘ��.:������ ��/C;6\���d���FEKe�����!HɌ!`���vX�5�oӉ���Yu�:Xq�T#��n��NN�,�eFI.o1h�E\��B00%��|�^�x�Ef�������t<�,l~m�fNmn	v�e����'�I�X��Lei�H�K�{�8����u���8$L1���7Fg�m�f��)%bHw ޹�y_'p_8zn�'�S$�ȏK�M3����5�2 V�;놐��d%�B�*����lc_n���}�D����(�樆$��+F���KwDA���*��K���W�K���^�������I;��*_��9��Cz�����M�'4:���S����hY�7^(t�g���Z��qx0ӷF�;͙h�#�X�鄪����\�0B�q���q^S$�5�U0f y��44\}�U��������#E8�iڬ8�5.8א�-:�a�c{�#闯��^�%���s�P�ٽ�S�(qFH؎�CT�*��[<�>6��{9�u�Ø�f<���"O�E�W�Oк/q}��4z���(>�&^t?<q\�U ���Sf}��%_c�Hf��/n)ksQMf�H�~��˔	��u�c�5xG�ʞ]TZTY�I�ɸHx\�t��p۞�W|6���#N
�%4g�v��V�+ҁ�ۍr�&E�/��AY)Z~/�x�����3��X���DlN-�頂3&'wY`��ļ�Б_�:���`V�o�����=�r�	a�MX�<�?�;��~�Y9|�� (�2Dѷ�!U����A�'�P�)��0"�i�u d��-��.�؎����2I`J��p6x ���c��8B���9c�<��~Ԩ��6�X���^0/�d9�a9�"���	3^����Wl"��K���#y�7��%�sqi1��S#���V�D�� �����oh�@�L*��Y��Ot�=xG�?�O#��UU@�[̌@�pS����E[q�Þ�`�lTnq��ќ�����;oy_e��e���	b�#�ݪ8�˭��b��Ͱ�2�FoP�CT1y�uG�jaq�\ߩ�wC�D���mvV��~X;�oഐi0�(GW�7򊌉�~�,�8>��0��}��������*��n�Yk��%}�7eӣ\!�2��4�������޹�S��&8��=;!���M��4q����8�Z겫2���
��=jsb�����X�$�xK�#�E�&������o2�.��g�h�7��hX^���;�L��Z�5Z�~��q����+|'F�c'��}/�G 9w�#��^��m��S������;�Ӵ�R�y���#���\#��'�ԧB���v]	s7M~��$�#-�:�!v��Y�����y��9�g�$B�v��cV~���KH�MĂ��X9���Z�_�ōd�oVQ�;V�M1��䗭��m��{<V2_K��Yj���yT%��b���צ���Qg"����=�a�}���4C�Z��H��������O��~�h=[5r\`:�:����`��T����/���`���5�ʏΠЙL�9P��@T��bJ���4i?ݢ����w�/�N��"a��U�"��W��L��<�4�������jD8.���CI��˴3�Y�8 �L�)ַ]�o�$B$"͘�ݤ�%�âIڨG�]��:w�'���1��5�X��>L.A��JE ƞ`F,9�p�ld(�:���\d�'�[H�]��7.CH\�Qم|� k��X��;t U+�q�^h+�AK$1ʹ�j�ߊ���n�F����A	�6���x2ϴ��#��H�D}��
R,#z���y��(pP��t�����������l�B*�`V�������b,<�76sm�9�����կѝ���ٗ��7�k"�sy`�!����
�yN�e��H��C2sz>�^�("�������,�o�h���@��N�>��=z]|�O�#�f}^m�MUu���ӷp�$�%���8��"�1jg\[���*�P�d�>>R����7���xr��ot�B�9����o� sN������Le4ps���՗P��D#A}Ê(9x5N��8��B��'��mq{_�x�����C�Ɠ�t�����ҁ����fH��M7x�z| OgF�C�U�S��f�٣����啨��cHN&����X�+@kG\^�*��o��Lԧ�,�{�űk�@hnKm�6�2�b"�nh>y��:QM�v�E�n3�n�r���z��=1�~��ޒK��cH�Z0����x��*���6u1�O�K1�u��r���7�VG��E$�I}M���n���=x���ۂ�� TX��"���:���%L!E��ԏ�y��c��!M�K�Bz����S��9t��.-�I����X�%���l��|�cRh��u�����5ǹ
��!�L�����FcXG���E�̦�$	����@ɡ�̙��4sl��5��������Q,����l�L�\4���?���������V(@a�1e�8���JPf���� �?W���K�[��4�g���RC��OƯ�X��J�$�E��]7��S0!�f\�9���Z*9�ۈ�Vz.$m�)��fO������v�q(�ІB�������Zf��Jn��\���2}%t��E�c)��H���Ѵ$���6a�,�O=�}>�[y+PpR���Q��8c�2���AW�ܠ��g�״ �r��~�*[�H��'7x`�'���x�J�=y�O4�@�XC&��a��e��K�����@f�0�B �l��vT�A�����L�
�G��d���>H�v��f��7u�2�ڑߙ�t�D=/��PLPθ�Htl���6H�V<6�D�к+���@N;<�I��\��VpC���b�W�x�c�������r�p;֨��62��8�!$FU�~�����6ϑ����$J���-&%��QX2t�Δ4�ԅ�zw��	5�/����A���1�]ꐕ1D��V�ُ}�}��Smq[r�ʡ�	N,�������T�d6Q<��w�Q�����ޠ���v�����!y׺�"1�)(?"<�)X箝�y���m��߆��RA�Gm#��O��o�3�Y�m	�'�ߞ�5�8�6_�d�[`8�Ц4��)Ő�).&��p�p�sm�������b�Am��>[h�o�M�˽�_��
&����8wbeF���w����a�)��!��hy�C����0&~[��:Che�2��9xz5џ�Sd��܈�?�<��G�R8�������v,���I�E.&ڰ-ۥ�|PN��4��� "�Z�%*��N8�?o�2���������/������]{-:�{1h)N	q\�6ժ}��gj�)+G���dO����رD�<�Ă%x�s̅�uK�[� ~�x�`�)g޸^v���以{Bv���W���{
bM�f����H=��VO<�?%F ��B�?����W�Л��X����7/ͧ�m�Ci�>�|ɒ길�[��&`��/�}� ��V�^�٤yұ	+�p!u:z|Y��
�@���<KN�L%��Q��a�Ty��/��5j;��w��*�b�$]�L�|<��zk��
57ٴ�=��8X���Ä�p���(�Щ��HZ��λGL���WxY���(xų:��~
���X���j���iI.|�?��M�� 6�Q�/J9z�8�rN��"��i��k���b�"z��,9 {ȟ�/cv3���=H���-���Ib=qu�$F�(���7͌,���Ҹちׅ�]�8�s��%�?0�`/���g�>���Hl�0t����cMk����$>%��i
���*��t	��x�7OVO�u�X�I7��o���:��"x�	~�j��W��Ŗ]?{����&Vk ��<�)u����X_ M�č�=A?��ؔ#=	<{�r�=f�_9��W��=�]��lch�<�R_U�벂ucg�ٹ�����V	`c��wBh���bʆm�`���,`����w��: �}E_��q�������6��F�c�C�.T���<��O�=�!)T���Y��\A�8 P1�����}�#�5��J-M(*��ecȧ�L�i*��#�zk
��C�*�����R�^��-����H;����1����;�c��ϐi�o��W@~�n��sT��!�����D 5 ��*D�9z�gն;Ý���w��D���9�'�'6��X��/�(\�IKb�D[�תr���q�D��'I���N�|8��H�c�J΢uP.k5-
B�]b�L�%�bEied\a�ݦq�S	���`7�A��g Gy���]g�U9�1r�\VAt3pғ%�h�tiڹy:�̗��*�~&�-C$��{�o��~��=!�����>����Ǻ�<��8AL�A5:럷���Ox���L,�2�h��x����xg���ݴH\�s��KxYZ�wdK�C��zV(`�V��[G�f�?��@�*�v���y;��Je���kޢ]�!��U�S�We��1�  �۽�b
;/8�W�3�&���RCQ_���B�X{�T��]�l��@|�]�u��.�G(g8�L�b�0������~"�-�x��u,���>�_"�� O�GV�m��+g�����)�Il����b�m��M�4�WR�=�/�;%�/J�����ȇԡ�d�������ʓ�Ҥ��E}�E	�p���lռ��6�rB8f&���7H���V���.69us��5-G��vcL-�+��tb�d2ͣ��=�� �Ш!E��SI�5�l>��
��RF�c㲏_H����� ����&[L��:�XMq}Z��^��T,���b�>���
lԟ����0�\W�7B���^�@����v�*��px����m��m�1�'-d��6Z`�Z}���Jg��s��ߎ��̴pO���/�Y�w��dy��[��J=����~�-��A!��$��{��L�A^O[���p�\��a�x���4:���m9C�I+�e��f�8Kt7�'j�j�
�z�cL�n]���W�s��o�'���嗖������\�_�w9��F]͜;󷰊W�k\�j���kE�W�X�+#�h}L�}.�ZhjF$DM���ԔO�6���J.��/U ��֙&-_T"kjԗ@+>Ǖ��J#�7tU�TM�X��c�MASk�~yl�|���n���Bdc鳿Gh�N�a�-���)Բ��4���M�Y�[��Е�����RD���L�A�z�K��<�x�FY2�M��&|(Ԇ���T�om����&Vg�,J���_��E���kӼ*�3y>��K>���
-ޭMc��H/eK�7�6��x�S�4�(��!�J����R��y�n����3�z��9�S�/t���	����K��u�W�V��}R��m��)1c���=�M�9۪���v�cQOw[�2]��o�Z*a�奄������%�?�"�2z4G>���Y�9�"��XN�W���9/���KM) :U3��i�ŀM�Y'8�>:����}��H��'V���8">H�)�̆BT��U�#�7����Q�U6PH~)R���T���>r�qZ1	�j7���DU�^����,�!a�Z��B�̕	��ZX�A�MH�"
�
��
��g���Se�Ϡ����h*���E �b���t*�I�Avc{���ҏ�;b6����ϖ�;0����v�U�d 9�p*D;����)�Y�`M(�|I��d���^Rkp��0Ɏ�=<$�O����M7T	����׳۹%��F�R��ٳ�R�ׁ�)��h�1l������-}��4����L�ڽ��pꎖ(i��\S�w>õg�@�7��Q����n�u`U����F7�������K��!���S�-/C�_@�i��%��
�NQ��l�8 ���������;;��:���S�~�S�p�H��f��l$��\�Bg��⺨-Ê���D:�#Z]\ܗ���~=ӈU��S��l������c�$�ǃ��ȫQ=��UR:�݊.Xz��ſt��Hլ�eC��,>�p�t�x��S�&�1��5v����a��hX������9�����V_T�^΃�>�����]�j6���x�%GvI�:�)�� =g��%��Ӣ�������t���G0�;���7��v�X��0J
5��-v�*��n"�淹����eP�z2��oy]?gT`�=O�_��#�88��C��챯�
�+"<������IC��A@v^��ȩO�n}~{����$��_\K�E���tJ�Iis$�8�N�Zi�/��6�ߗS� ��\����/c)AeS�4'P�B+
��Q�sE����BF���%dz�C��.v"���� ������ƹ���Y���x�s����� ��{>g�a��>l�VaV���������\6GB뵄�w8�w�4�y���Ӯ���CT��/�z'���v�Yp�A�	=�Aȑ�f� �㳩��.���(r'B@$0��Eg���IV*�GDa��q�0�g��t�gLA%,޺�ߎ���y���6[?;��r��)<��5�^L�9.��M]h��L��F��Y���$Y"�J@��!���Gn/2�����vahY,|�$��/fe-ъ
��&�:���c&Aɥ02v=;9	ڏq��L����~�R����w$T*J�nx;'��i��m����N����p��G��gu�ˈ����6��^Bb�e��������T9�|�h����9�:�=@M�]<k��?�G�;p�
S&�5)߰��Zj���;��>6�{*�_(�7h�`�e�̦���D��;������h�Di}����P��dR<it�F�����W�?�rtJ�ƒL�[�ɧ r���~ෝA�`��D�0�����]Lܥz�6�h��<�E�-��y�<�cubg������6���� ��Q���R�D��,�QxnQu�����($�2�W� D08%�pھ����R� �L��6�*;�)����,B`ZQ!�?ㆶ��IK�3���P
��[}
��/��~�k��[����m���i��Б���p�ö��74(�d!�N��ƴ�#�0�69�_���Rב�-�2���_����X	�*3Z'K|d���块�����<���7ƥ�l��R)"�o?� m�[����d.�l�7C�IQ��G���H���������nB�����ٙM�.츙t����Akv�K爤�5��=����0XJ�R�R�^.�Js�=�PO^b��Rꀓ>��}j�^�rs8��4�;"�#"��2�w�{F:K����$^?�ee�:����6��ka�W&�({�8,�%\+Q��(�vu*�����ƈqL���ҿ�KL9��T�R<�������� L.v��K�ЦOՂfw��4�r7+��!ۑ	0���r��Tb�x��,V���)�e��Wg��ޫ�3���*\��-�d��}u����������0�&Dtb���"�+�lL@s>�6}x�Ŕ@�������]ݠB��M�c��E��D�\� ���l��b�P����v�Y�-�"����8m(��н����z/2�.J��2jme߼�
 ۙ�I��iY������^P�帗�Ø>l\�oj��7�/@�Cf�V��� Y��u�>o����)h�9>�2ӊ!2�d��
Ru=9�%��e) U����xu��UeDq�;s�X
�
��П���!�5o�f����!�	�i��}���cv��;d��oI6|��R6���k�5aF� �Ӥl��j��L=��l�v�%�V+��N���1^��[<I�C�C�W�ǋ'�R����AP�r�\��Kg�R��=����I.�z��`(�b0�8L�t ��~��UU{X ����HA��nv*.h9�㱈��pTb�ۜ\�1�
U��uJ��-σn0v����c��8UR��	
u���2������2�eǽ��y���vҎ�z�����]�ʥc��ߌ�Ԋ|�1662���S���b��S��$�Ǒ��r��AG���2(�j>	Xf&�<��ٷ�T���3}��I�e?T+94�{�%ܽ�ޥD��/�	i����o��B�Ɛd�*Ft�&�Z���AN�S9��o��̟~�1;�w�YEm�ژ�h�D��I���V����*�9���^Q��7M'�6�o�^�U�k�&�CbەΗb�:ؘ�Z�/��p�q���A���2���{0'xv����.:���p(�������x�~�7�W���LHǪ��ꎁ=Iv����rbe����h���4S�;���E�V
^���PAaA��h?�H���>�&���/����}�'Ń[�9�$�p��G��f��]  �^&���t���������P,`EU�`�3b�A�?	Ʋ>�%�,�xВ�J��՟.��V�����jZ~{�����Ҷ-:��-�x��Y^rE��򝄦��?�f}�r�z���)N`��s��ZGLE�:[����U�&H�P~_���}�=��W" H>��D�G��*O#;EVSxO<1��;��)A�/��E���o��`�&M��q���w�SU?�+_f����$���Q�9hW�����ҡ@��OE�΅s5��MW@F��^n�J$���o�B�r��i��1��y�Ƭ��0�9Vr.s-P��f�3�T�N�w͋�S��Q������yE
۹�r�{���ɱ���j�gZ�:�%���un|�z��#����Q`.s~�~�gdhn$bn"V�c��@N�d��؟:�m�!2,���7ґ����l�د�~:i-�\�c���騼u����0�C� �,w���H��MLo��2�@��fW�RV\��U�v�e�Ն`c��y��9��hWdti-����\�Z:����� '���V����N�şWTV���T���u1����<cv����g�\����=��[%���z��� ��fz<)�l�#�;JP{Z���i ���z���`jA��r����]�]�$�� �t=zP����!?�ʢ��-�����`��~��"�����>�C#Q?����-)�?�6��0���G���S��%��%J*�A�	u+���Sw�Z1��e�!Ã������I���d-�%�Θ���I��+Ohe[^|&�T#�]<�?�0#�=a����c&�<-�_�	��Y���d�L8�����p*�M�x�(����`ަ+��Ls���<U���!�r�ޯ�k��)lL֓��ן�X�}�׍�G�˟��.}<�{L�#���=�9��Q�Q���9�=�,��7[���m�|�2=����d�c�N)�p1��~���M�Ǩ����Unf�7�0��>ڽ��/{�s�fw۟��BE:�Km��c4�BNV��AMox0���eΟ\���.��g"<-v++�T�>�%���1;fe[��Q��2�՟A.{��={�IH{릟�O`L�G�/h�)�1�7��n=~��He�,�.]Ee-�H٠��:��2�%[����We��4�@n%�l�F�_;I�)�漡��N#� �������\�]瑅=:K�l�c�ɯr���&��}���Q@�����fE���}���Y��f0�{h��I��Lm��+޷�����+=؞1��*��{e�n��/6��^��IH���-툨�F���S�����1��2�tn�.c#�%��h�s���36�������<���=Tb�"�0��8�|Ҭ���?�lI���-�PI�t*��d��."^�uI ����`r [-���
�Цs�����f��~�P$4����<C��ؒ���K�?�_C��a� �VrX��U{M@L(T,�vi�J�Gc�^8��L�J�����hV,%���5��m���t�^�##�79�R�&H����B`�1�Ngpǣ�e�'"�Qq�Z�_|`�v�A/d�5h��Zub����k�l�ie�H0��9]Ġ�`,��!:b�w�Fx1%A��VD�j�w�Զ�Y�W2ī��������Yl��Z�ڂ
7Q�hj%G�f�Τ�D��@��I�����l������J�l��,��e��}����μ�-ư�Q��	��9WʟA�n�]���V;<���R�������9����� �-�?��t���ɍ�E�	���3Z)=b�d�@B,�{�E�������ݽ��L�Y�)�(�>��^��R��ImIo���*B���GS+E�|���K��h�����K�>~~����]V8	����(�`a��Gߖ�%S����T-�������C��d�6O�}�šh8��e5�c1B9��ZL�"��,�^8�7f����ڇ���6۞�@rStJa��%��^���胙���/{ 品_Ŀ<%�T��&�� ��7�=�n̾������]�ڙ�Y��VԔb�7�г��R��ܯ�)n��RNt��w�q9�8���uS��	6�0gM�U5"Y�[�E<{re��[�d~��D%�O��u��bp�>(Ҏ$�g�F��:�3oVο�>�󝧮�T���i�A�D�z�0Ԁ�t������=\�8!mʲ|ʙ+��K��'8p
c>/_�"�� -��OA��L�#[1�����&�=B*���P�"m]~5`,��?l�.cW�˧�BZ�d�FV�X�}���_`��F�x!�˱{;�n�'���}̇��̶���>�Rof�XZOqį��ZLˡ �QZ,��6W�F�c�N��I����	{X>eRR��$�4�m��7���&6/��Mޙ?����ƟC�h{0c�%tk���ˋ�����;)]�P/�����Byl��f�#<rtpk� ��Q^�Z��%��
��UX�F6���?�hj�1�6�qt��O�;��E����ZTѷ9�l�Fպ>e������K�ARߚ��̸�4Oh��W�AQR�����F+�Y2��,5��T�k�N�8�%�N���ݼ0��V�ӥ_u^�?~�Д�=��%8����;�j�dWq+�ܞ�����~q�-���z,�7{N�>R[�M��F�K�БN���^��Q��B>C�F����+CJ��k)�f�%��a�Z��醉5Vn۬/��"�*�3]>G�%q����ܬ�q|<��]�>�Wy��4�Ku���4�yR�oc� +p���C�
vK��],s ��7�?S�z<lfS�o<�R��Q�&�:�� �;,.��� Y=�]�Vw�)�%�(���wP�IG�F
�e�6V�8��9���o(�{���u�~jjHKD~@Qc��
�����9/���#������Y�Y����ge����L�F��:�z�L�w���˛��|����38�?�ޟN�n�Nz�.���П�n���E'���N-��Uc��E�MR�
�e��������r{ # kp���cM Y�}��%R�.���]��Ȏ�<��՗g{,�`�����nベ���U\~VE~�+�
�ϙ�2���f|-J]�$�K�b����h<4'��#�a�nϗ凫�}�}���gK���T��{�}�"�f�ٕ��Aŭ�0�{�Y��_�c탤�k
{Q� �8j�����2B�Y<���0%��|w�+��ӹ"yf���&��F�|�G���:��1��TX���ZD�V�aR���}��m] �`�B�l�(��MJ j�� �����u�c���S�Lϴ��5�����(t(~�ڋo���ԭbR�fO6�K`��5Sj�J8��[�D����[��-E�������"��0��w�-a�k�֧U��閭_���BT��7����$�Q��{m1N�K�X1�e��<���������U79}��A��{�ٰg�sX���N�p���iWc��L}B�}{J�UL�V7��8�r�����w_|����>1Y��%AV��qXKS��$V��[�z>I�p}��)D�Vw��x+��'�7E	
��A4�����4���g2���SaY��1eY� 2:s�~��(�X߼}\��_P�`q͔�3V>K�1�!����1�%�p|�N=~J�?PP��;��$��1��o��Z�Bo�Q���4j�9���ݘt��s��Gt1�e��pگBq�%K�	>D�`�N˱��n�N�˘K2	���p�Ơ|2�@��	���6��n�E2�\������ދ��9.��d��46�!f���,��:�x��g5�A�=˶�����§MU'�
bB��F8���p#!����l�y!�ᾣ����Z��ޚ����2�G�j*XO!��d�2�-�e۸[���g�!f��/�����2.�e;���ō?�Ue���"WW�d	Y�L��=��79Wڟ
����RW�6��Zz��?�1�`fR�C%t���h;F���$5KS-�d����Ձ
jrR&�����Yz�5���@z�7�YF`L{�B>'�Դ!��C��K��O.���A+t��^���L|�u�p����P�-�s������!�Lysө� �`�)u臔��}?o_��.k���BA<{�B����ww�nG��тP:Xʐ�-Al�h�3�/4��&���a~�s
�T��)0�-gc�3�tx/���&N�*7v���F w�y�t6a�#ҴlY	?�w�0i�O��e$^Lh2�E�)��G���g���6��eK�/��\о�Zp=G��fqf��S�h<k�SI}���qr���nFmAW/���JY}s�~��;�>׉�'��(]������1� �yn��ٟ��:�|*4���YM��=���&�#��b1�Pė��.����ț�ϸ�0�����2�
���
O�)�N���\.a+T��A���!���L7jpvد�;�@_yO$â��(���1�*����y�/�����S������˥jY͔����:�4�_����h�G�-eb����+��,`��eǀ��p��٣�]���濸)-��S��/0&�f� �e��L���Co�pW�z�>��:��V[�ڒNO�oʼj��幨E��,a�Q�aj��������Gz���N���s���R��iw�B��>%�ٕ:����H�ȹ�X\޾Ԉr:�ȨD���f��|{���|,٪'{C]g_k��=�wؚ�f߹��\���Y���p�ŤTO�P?0I��gH>�h!�	K��^W����t�>5T��w����Ō'O)Y���Ltz?�ҫ �Gg�����j�hH�*T���m�����D��L�R��u\Ҙ.=���T_( :=�Ro����KGR�@�ʥ ��@���Y�E;SM)��hb�
	?j�ճ[Ń��I��4q�
�̒��ʤ�Y��Խ�*�hءNE��h����U�+�0 �7
�jw	��g�i=-b��p���u5Y8:��y~���rL��j��G�o��m���SR�s�T˄j�$�M�Jy*�%}��y�I��[�5c��& ݝ�V�?��[E�Т��+O��V��{�x�o�	���C!�&B �t� �Y(9�Ѭ��@�������-y�;�| X��8lΩg�E4Z�`�s[{��`���a'
�5���H�kT���_a0~p�>�����R�ǖU�����U��z:Se끣�A�`T(�i�	3s�ܻEY�^�؛���1��=`��Y��rL���o]��s��߿{�xͭ��z���D֢�ϝ\ƨsou;[!���W���r)��\ .!�����N ߰�Y~��z�z <奭-7e��]�g�r7dh�xp�)�����)Ivߟk��eq��ßL�x��l�6F�|����M�v.T�a߬�ֆ��YB�J9�t>j�?�9�$�B	x&��� ��\��fke�(O�����!�[#`)�~eS�>b�̃;օ@��g94R�'v!I���hE����"�b���̯���09�����#�x������v}K7�KvsR�Q�Rʛ�w��q��b#_�����@ޱ��*S���'�l2_�U�X�(a��I���v�|r�9�X��*3g�	�n�:H�v|��r+�yФ?z��Ӽ<9���Kw��#�[K��㹔��iD0��FL3��.�6۝�b��kl���� O�3j[mAq\a����:oD6#y���J��P�\3�ۆ�2�M�;S������ I=M���`��K�H��W���.jϡ�ud���Yr{~�rr��z3C�{Z���1 �l�B<��� ����oZ���ܖ�i��M��G����~��	��I'��x���B��T�Lo��}`��,<��͓�I������(���o�?�	�9=W�;o���� �w���� ���Λ��<���[�נ��.��Ĳ���я���[�z�i���Y��wG�w�Y��j��D��AdUy=��,�usl3�1a}t��|�Eli��(�j������ӳ��Ȗ\3T�f��`�;LJsl i>�D�5�h�g�8vW���p�OBeح?R*s��+L�r>K}
D�ي�����Ȓ[�������n���K���%�8F�_�X���c�q�y��׎�xz,�3�|�DV��]8A\U�Z����7O�� ��{�r��hR~N
��@xr�>�+��	lD)`�>����D��(�����)�y:��ڮ6べ��cS��K�\���a��UK��i˦F0'�,�NT]
>2�'�KQE�V�,%Gu�O�Uto]a��8�a��:����S��0$���`��R�Q#_�Ƀ�o'��
h�]i{s�&��ے��D�ߞ����o\�ѥ��A\G"���s9�uM��PBJ��6�G |�:�8<Q�OC2J5�cN=�.T�ꎕ)˘�����!2�Qm�5Js��|�����/���@H9�����Rz��0D��貼�@� ��W�A/I_$�	M��g,`�C��_is�lS�Ŕ|���Ը��x��lcO��@�SïtM��'��NA7BY��*,�
 L��M�#��߂$��)�B��z�û2�o�W{z�?� ����v��QU,.��~��4̍� ,�aV��:�_
8�3/��Hm��ݶ�\���e�}a��h�~�ÎVT(�=��HI���&�́IO���7E��&�~�4��������!Jt;�<iQ�Z�󎹸����)��J3�\�];�Գ�@+��M(@O�#��7H��J�?%*�E��__E���M��̏=9�P,ۚ��������m�V*��<9>eBo�5
jۼ�3]��j�|P���(��7�U��b�3��Τ�����	�a>���5&����1��bCg=���-)�m�;��;�1���w��60|��d%�~���Psn��J�c�b�Uk������:&��Ao��u*�6�P��v��}I�E� k&3hy+x ���[�����pO�s����>:׵5�?�Ǻ��`���\�p�)s/,�L�p�'7�'�R��ʐ�m���R�N�{��-��!Ȅ��3�>,����x�d� �\�z>Q�"~�P.��`WN��랬�������#	�Cl�y���p��B�̼��M��Y�xr��}%!ؽ��������.{հ=�nK�P��^�cn�܁4�2H\�E�+�����~�*US��9��?��b��|$8��xC��NRE�4!���Up�h�����PO���Nź���6�7����f3
a�3}����U����l;0Ƽ�K09�f�8���O�h��%.��֯����^�J��[6��8d������?F8#)���*`��dq.7���չ�	`�g.�N����< �@#@�h�-W,o�	�ǷW�T�%��c:�a�Bb�&�%u@�X4a���1:��GW<t���%9�.`�����ZS�R�,1��y]����ˤ��B����P�+�h?U�tv�$ヵ�i��J�����d�Es�
�9u���	��H���	E����zJ�K]8�xR��4N�񃤄@�T����&��xL�yn^?ǀ�[�3|����w)B�M��p�ڧtҥfI���Q��Y|�����ՕCm&��6����%��Vry�\�K�~t��& �}c}s�[�zo�P�� ��v���8�>��%�� �!(>JXK����+�R[xv�C�K��s����J��u�������D`�N�u��o�Z>K-8�˼H�?dˊ�����-ڲ7n��*�0]/@�;����Qf�r��%R"�n�<
��A9����u�\�2�%�j���$70a������M�yx����~����p���#y��1��[�(�ݜ��8�E�ANIƵ|��vLz=��M����<O�o�O]��<�@v��u%���=��P ��z�&���]�-3��s7��_?3�]�G,6�LB2�'�1=���ƒ���bkd�^�WO|db��#�Ǚ�3H�C�[��3�c'�:m2���> �R�s@��D���6a���R��{��_z+.���'�w�	=�E�����h��zBF���7x�-I���oVI�������8H�3(�Y�����}�▊v<¥Oba���iNM>?t��,�~�W�a��k���g�Q0�R����U��qG��6��;��}��;
ѱ�%�y�9��x�kɾ�����s�K��Hv�*쟡�k�$�Qu��̷6� 2��!Tn}�p�,�C ���-Ts����//�#�Kb5j-��U��*� ?�'tr�sO�]c4y������n�]��It,9ʼ��Ł�(�ۧ�C��Y�!oį۞+=^�;y��C,�U@�h�}�<R��sS�|��]Å��s�����Ho���1pB,����%�@�h$�������+������X?:)�� �W~v���x&������k	
q<��F�G߾�XD���g[��Ѽ1Ƈ-�9h�=�R�ߺ���9�%�پ�����n��w-�W�9���A��@�S}8I�����~��H������r��� ���#����!E���b�u:�OBvsr7�)6��[΂���q�W����/��;}�7L���FkPO4���p�r��8&ۀ� ڜ�.=�[�G�!�������42h�lW�x�?�����1�doQ���Ei��F{�z�ǵՑ���A'��/����t@�phM|�)�n�G4�8�A.�>p|�������'�%� n��[f�0�ۯ�tH���}��~����X|�������A~�;].�o*����D�Ā��S �p�}6��(��X�P#��fΛ6�r�[_TX����z��I�`n��ْo���$B�3�0x(��n�sr�f�'�wJ�M.���ec��\d��gtv�ng�\
X�}\`:E�7.��^��w��	���Ne�H%Ѯ�*����=!��BN�fPï���\������>+�_s��5�)~��M^�$��3��#�u�$��i�dfN!�,���:�}��@n�@�]LFzL����۫�����Rgkf-6��i�O��{`�=?+�0��u�Y���_����!d��Ap2ʓ��9����bY-����8�z�pW)5/���%s�i��"qv��2\�<� [�qԛ��X�H�����g�&�>�:7R!b�V�r�^%Q��^��0��oĔ�����#���+m�t�z��]-2��X��Á&�x�mV[q�ͨ���7��Z�~��B;8݈�;�?�į�?��Ґ�F�>��U~L��R�4>�V��{��hG[Qҍ-)نQ�d�-���9��< >���&�K�v������u��t�Lj#�V�R�*?ݯr��L�5rUF��TM7�d���w���hJ��'C�lq���+�A~��M3�Ͼ-���L�Lx;2���T����?qS����ܳ�*Cl�[�L͔-n��,��ߍ����jr��>.z���}{u\4:�S|��d��M��"���:�NVD�Fa:��dսV��Ƶh��?!����i��[�H����!H?��������.t��{���w'�,�nJ�5eӰ�5.Uܳz��#��!^�'V�&oo���e��[��ˮ��`z2l��9�� /���F�dZ���9�s�|��Nh��g�<:i
���5�ӓ��H��a/��S�Ԉ(A����h]�|(1�RۀݐsZ��ѹ��Vc�>�J�c�$�=��
�g=�E+)"�׾̆��j��t���Z��3���Y��ĞnА��jֆ�V��#�"�aQ_��(&�P�ںG"�8�D����}d�g�B3��1a����8�>�Xe-�����x�Pd�9��8"P��
����uuY���掷lZ9Ra�[kǒy�@�[}!g�@!�pR<h��1�>�Ϥ��
��cU|���m\�;� ]V��b��{z�[�t��ۘύ�{���ް>i��bj�7�#:�5���S�C�j&3�G��_]�XcA�駇�럎.|�����r �1�X�Ŧ��l��d�O��s�[���U�8�?�XD���������
jއ]`z���	���& ��,!�-*�i�O�W��?+�x�aYF�D�[l���O����1A�a��sZso��.p��'HHJ�q~��zC������Bdl�AC�����t}y�U=	�&�_2��Z��cװ&Z�N�/�"D,�&k�R �cnt�&b�µj�u �u�S���s{�f<�A��c�p�'��G��dT�XrYB�@\x�rP��\7�k�s�2!~H�����@���q�;�K�:e�{�*j.p�xre�;�= 3����B9E���uwn�g�� �MW7�,}�5GJ�u���<%�7�5�dl_:�'זc����ǻm?1=V�d�s���:/����j�����<q�U[��Ûԍ�2�Q�O�&���Gܿ�������b��4�@���k�6��6��DZ{�EU}�\IH����0:r	��.t��C~^+[,ޜ;&��;�D��'�a6�m�w��
��6����ܰ��s��t��N����w�3�W���&��?2�������5���#e���(�V�%p��ʟ��f� ��u�:W��^�9��q�f�.O�Q��Y��	٘��"x��N��2���.�;�t�;�Rv�3���{r�YF�����U��U�>$�0WL�mkXSK����RK��2��H����z��*�Io(K]�b��sL؎'	2d/�@�5��G� �#�F69m"��v��Ɣ��~���.^�N�A���C��'���s��|��b	�#����p/��y��;��s��c�\K���K�{���r�C�����
�LTà0���Y�� �-�7<5I��އ+�kw+�c�0X�خ	±��.�}C�����UDXc�.�C��� ���F��EV�7_�u$y.�r�Py_��)�q�vaί}:��h�l?v�P���4�A�næxw��dS�Q�J�}�h��c�BۿM1�E��V�:�G�Wp�I�r`s��G��Sh�y;|�9��<��If�D`:Mns���B�,0��EbPY;)����]� =c��b�䁴jC��i�����|�� ؽ���u޽�����R�0��[�0ା��2Nc����Y�,������bZ2 U���bw���@��m��J�C�2�{��)	�sJ-|��ߥD� C낇��q��sO�)�7�$�=��X��)C7X�F���W>e�`�����w[u�t.�����ݲ�FL�ey���=�>٨5�jZoc.��o���5v��`��-mޯ��<���p	�n��؆K��Hݹ6�������Y���ۂg& FYv���q���o�����g^�]!�~/Ҍ��k�(�I-��;����oJ�6�12�]���ȧ� �9�ۚ�����lٚ~��\���2J�n�w����G��n<�m���.�l.�O��"���bF������"�<-.��;l�*�Y.W�-�{=�\���Y84ŭ��V�R7��L�� Q~�_��7i��xO:1�ɮ�'�*y'B���ê�nz��C�Ы-VM���#����T]跮�fâ��1�i?�s��o�Dd�5wpt�Xm�8���,�e����~�/��{E%��}v}_.�]c��$��g�?�Չ����+��<��:�.	�Qp�α�#]7Q�X�E��`�`�l����QK�dL}夦��w��FQ�EY�`|���l���T�G����G�@���,2c��gNmg5E�1Q�p�����n��f�S�]'����\!�T�OG{89O�+<�!� �8����_�M���Hlٻ^���!�@N�Ь~��D��:6B�zq/}h;x��X*�\jam�a�=,���֎�����/f�*~ja�.��bI˨`��ٲ:���.D��/[�����G��Ki����˛QP0�
���3#�އE%Y��!o�}�mϳN.�4&��uQ����"_\/P�oJŹ�bpEE&eR�	�x�(��Ӻ��04E-z��D��Ԝ�TM��ս٣�ش�@�[XzV �L�F!d����Cɻv�]ƙ����|��鮰˃oK���=�<H�d��?��dW��p���UB�P#^�g*r�'f�KDο ��{O�a�ָ�An���X�"��v��;C��*{�!)��S�������x.�Nؑ�1�k���ȟ�*�&v"Ѣu�u�F����v��!���qj�ܙ�b都�lR�l�=1F����]�?�D�J*
�%w'N��5}Ѽ�	�ۮ%9`��������"p��:��N�_d��dy�0i�H#(��"�_���׮�{��)8S�9��e���{��#T�@�ꅒ*15�K	�O��׾�rK�_��&N+^��i���)<�AYn}B����;�GO:��f��`�Ѹ��)׷����!�5/㣌_O�݋b����saa���?Cj����dM��Z����Z���#����;ʖ��r���7Đ�Ҭ���s�Z�u����.�jL&��l�$Y����9�K� �>4e�d�� C�ʵ�EΜ�yB����+Av��ª~&|�ݔu���H�t�)S��.�7�h�C�	�fg�ג���3��X{��9� ��.���0�ߘQ�p�II(�k{p���)�Gt���o���N��L~0�!#`W������� N߷+�Lj8%��}�z�	f7��ǣ%�f�Z�u�n����s�d�@n�7���T�(k�)�Q��jF8�LHX0�k��f�=\f� �^C��6�u��w�d%﯐|���<�!�X��/�z�}YQ�(�?���w2��ȩ?P�	�����ίo0��pЊ�V�x��<R�1��f�9�N��:4�)�>b��kaoA7oa�w�P��#�\�I��(��V~�x���R}]^��_�a�yLI� �&O6��P��s�]:g�X�i |7�\iBx�3�C:���\m��+yu��K$�ڣ��a��$�t��Q�QVA��3ȟaV���J>k���d�	.\��ļg&�r_��ˌ`Ѐ�i=�ʜӢ\�<D��(\s���cln���Z^l�Jbp�����n2�����͌�Zqm<���y��g����.h�e��`B�P�W*kl�^�g�n#�1�+J�}� ,;?#ԻL�36e1��d�H踂�]�P�o�L򽚻��!f�m?�W��I�GՋ��<�1\4C"��,>¤6g�J�_;bH�vk� �����,!����*��=����o��X>D���ǵ���D7���"�^,l��&m���F)�lk�Eo�3/��D���}���f=�UM�O�R�-���'�s�o�J�»�YR��"���(?�`��(>9��O�D��Î����]���XZ�.7���V.J�T|ut_M�V^ƭ�{[ |�l�-��zJ_K�
��b��ZD>쫊������U*���Uq�%"9��w��M�IK}M����"�,�/ژ��:c�U��� ����u+�n^b�����b�߫�.ş����4a�ǲ���@uٌ�=.8�=���߰���v_�& |� <�s�τ	��:���7z�o�{���t�Lk �(��Fta�8�GŃ;�F�^��3��.�,/�{�p���Ȫv8`�h�}Re��gC���5��p�����{7�ƾ1B!��
��a/��b�%Y�n�tη����˼� ���4O���d����&3�`{��[P����qO�O����)Y������z����%�8���9��9)(�C�_���aK}WE��Vr��B\������>v�7B��ނ���%ץc77돈�ۣLU�ne,�F��o�ݪ��Ѓ)-1Du� �>�
�����,-Y�qU��$��UW���C�ռA��r�UIə?�w�"�8�x��m�p�aԞ�� �C�!��%��/�X����y�ܿ�4tE��g�:֐�78��G�h��m�ɨ�J*W���J|�ڵ�3J����b�5��Qԁ�
���=�y�j��^R�T>�
�sO�显#�#�����O;�ЇnS�HڪLӮI�����l|�N�g���6&���<<������]�����u.u�B6����ʡv�bC���x�@�S)�%?�������Z��em�`�4�u������J|�ӊ��(tŸ;nL(�dX�xZ�d%jk�ұ dڒc��c�W�FC��T���O>d(qjV���eS�*&{W���C�1dG�e҂ ޽�+��i�)�ě���0ɭ�iO�p��l�9q�_��@.�iF���O�����>�D
t���B��NC�P�v9�:p�S_���ۚtn�H�eq�l��儀�D�.m�����Q�I`�0-Z{�����M�	�gDk� ���/�Jva��+M��X�mtx�����#'����*����U�ue�q���T &5G�C���|�r����D@l	LP�~�鲨�7�떪c@�:#�g��e�j�"?�N��-�L�(B���'�հކF,����Y�팲r��Y���ǈ��fu���>x�2�9�M��G��berYL������F������[�P��;D?�2\���
�Θ)�IbwH����l4������ɓ!k齧ɣ�R��(����ye��u�f"�⮿0_����@Х�wc�Z����r��D��u�co�N�~�����Mbe~^�������l�&�颿�.!�����I�DE�h�z�\�GCy�2+������~HL���^j{������^e5�dD^3�/x�	������<>F5�kjC�_��M�i�61���5��l
���qO_͑:n\���t8hil��>]��ĉ.��9��Q�n'@E��@�DYc� ��+�;L���ltG(5TN�4i|�YD�ٌ�6�$�*N���h(y��蹂G~���,M����;	�F	BT�r@�Z�գ�00`\��H\��.%�iQ��)l
��=�:��N��V�ѱ��S��S���ۂ֩܇�e��)�o��K�,9�Z�|���\ o�-�K��ꆂbO7C��妃��U'�>BF
-ez,�^��H�C���������3K�f�b�7��M�������o�e}1vy]���������}�-̇B`<�Q�?���ch0�!?��p/������� A��!
�������]Ǘ�i���_��WJ����9.>j�!���*��6lk�VO3��V��(�u񫜨��k�*��HN�|J+�]����=��������#[)?X�\�,�#$�Ǟޥ?�kg��tn�/x��H���:ð�Ҟ�KmTנVZВF4y��Yh��R����׳��uz�k�K�OC�'s���V����e��aD��wc��R�"�e|��:%���H3����dIoo!w�Wʒ�U�Qg�\��W�Vӵri�Ʋو���łW��B����`FXl <&�)�w��jcU��	�݄�꾎�-)
�b'��0���m��R����h�n�+8'����MM7��%�sG�$�~}�+ߦn��w6�`z��'�<d�Ն�V2ot�n�fx��FhЕ���̖M �#_io�鎆Zk4|}pżunV\,M;�<���9�V[A��҂E7 C^LD��{vĻ�Xa^��j')�D6��)Հg\���>�k��k�AEj_3΂V�)���ɖ���y����a?�w�9�:�{_z�2 }���>/�0OPW9k!t��M�q����ͻȄ�@َo�m�u�
��� ��O�lzœ�&��d���c�~�-J���������
��o0�t�z����O=x��+�;��C�KR�ᐘ0`�>M��Bؔ?^n�������X��Y`�Ŕ�m=�*$�W�Î�;S'D_��=�PS�㼕;M�m�I��I�$�J������cg����y`�~T�i1���nHl�I�/�����"1Sa�CR�X�1���K2�Y�un�I�,�K�='�R��P1.c<�Q�Lg8ٍ�m��dRKE��bA�sՊN��,N�y�&���2����!毺Rщܞ5m�s�܂�D�2�[��0�p��⮒���Ă��6�L��L��'�Q��8p����hq�(�1 ���ݟL56���X�'K�)l�Z�gZ�pj���s	����G��e��������q�ox��"�X.���]�0�a|2n��ɬ�2�,��?ùU[T�6�r�E#�@���6]	E�=�����-��J��m<s��l%��ˊ�QP?͒� �h�e̡���N�W�z��N,0���+������!�F��Y�&e���g��}��H��U�����8B�&;�~��z[s:F��l�8�E���-�`:���8GP���KN���m�Hzlʲd�稧�\���{����,��ƪ|C^ţL{r�����[:����ǆ4g�]�:|JF ������[Z�3��%p�΍&�ę?�:G%Q��9���g"��S��` �I{�y|���ΥYB��F"��̂�o�b~|iWo�%9~�j�w9�1�n߄�\�]�r��/VQH�у be�Ö�-��4]�|�~І�0h���Vʇ�L+s��ҷD����Ȗ|��Zφ�+��U���୘����d��qZ��u�
�m����*�j��^Q* ���C�����~��nm"u���p`��r���)��\8+^n驶�U'ҏ�]�-ה�}����W��w�5v������0Wp`�g�2��[HB����zh���6��+�u�N��v�r8�~:V��6�Q��jc����Z� �����Ɍ7�>W !�U/{����o{�7c���G~W�YVl�qv�=.�K9YW�Wc��	>+4��;<���͸�1�_�r@����G��t��b�^�9���և�������*���t/R��wbih�PD�[u�JB�0��zq�Q��/뛟��%�9�t���K+J�,��J(1�
4���Q�G_�5�e軫1�qϭ7���+W��,�Q�b'˜c��d� :�)"�csʙp20�̑���@�y�d�;ʫ5�RL�܍V��\�d�*���hB����~�J\�E
{3F�&�#+殝َ��z�7�p�x��朗^�A��V7��EH�'er�����Ȕ�> �t*�й�NtD���f�]v�&��y/Ңһ	~�'�hM�7�Y�Φ���ç���甹���RU��\Y�$W�aΰ:�'���f�R�k0�_c/>K���O�y��!��4�WȤ��)_�j����^_H�I�_mf>�͠?�ӹ�j7SV�b�JPYRA`2fX5��%}Ǐ��_y�3_^Ԉ���%u����m����{��HSR��=m���ʃ�'2�j�� z������9.��C���.�&o����i�GNp��E)0��_��:����+A�$ѽ�s�/�� ��`$+��}6a�y\Q�mW&D;��zh%��?�bJ��-N�T���J���@�
I�$D���f]Mq��)�~���/r�&�?z�2՝/�����λ�`È���@_{x�?Ĩ��uT(�:8E�47n��*& g[�w̴�����}z��yi��@ v(����1�:�pH(o,HC`ի����F����'׵�J�I�u��˯Cy�|M�b����
;��SHA��RqjX��]�!</�,X��Ho���XW@�����n�І�	F�Ũ��p����	t���(�,�ĕ�ĳ;����b?�����-�@�i!,���s����NV���]�/G^�B���xrh~�	�����hV���t}#�"�5�?�.΋��<��K1��`˄�+q�^�)-�|��M�$j�]_���]�p\���V�~�M�L����d�����ד��D���ɖ�k�9f�1*�>T�D$�Ff��1b�1 �+�z��E��{�^*p�����&�Z�������<>	Tt��)����3oJ��-��?��F�JT\ޤ����9,�S��;��q��@Rƹ���v�<ߏL���h��L!��
H�>J8�rJ��8$��u*���ª#�m%Y�q�`qt��j�j7U�U�5��6|�
����E�"�p�,Ĵ�â��.F���!���1��ǝA�)
��������8��K˧��i�s�B\#�x3Qa�aÔz����AS��F] ��j��9�e\�Zk����s0�K[UZƃ�V�j]�Uy��U����������ك\���X�y����>0_�|���Y�"/ׅ|���挴���P �#���&H�s� Ҕ�Pc%9�8	2y�U�>�
X�$7Tͺqǫy[se�I��`��	��{mo�d"�څQ	~n��I��ǐ�_N�	U����_�9���&��pȃ�{*z�¤@�8��;��/�X$�
ry�cy��h��p��V�X]��؜ܬ���fOn}�yxJ�gRl��N��˻�����|+���q�g���3N�+�s`�Z���eM����ɶ��T:�'�C�3�o �.�^���{Xzҷ|�[Q ��(���G'`�Ɖ��w8���T�T� ;}W�RcH
1Y@o7�F�>�Ah�9l�T�4�����b�n鎘�y�%����Yz�%K=$�좬 ��]�����������>��Ҋ{Y��Պ�-X����Õ��˱=2(�>�����5��_x���H/P�N�=��w5|���(2�0��9������xn�ڊB�Y�O�n�����q���k-��w#x�|�ې��}����S������q������$�5���j�+q�sO�D�Py��PH�ї�y>�ʴ��v\۹��3�	��u��:���:!�,/+:�ƕ5Ҷ��ʜ��=�%��R,~�kl�˴qa^8��Uc�bĔ?v����Jd�=�(�A4#`��Ӆ����|�;�����̧ƾ�|$0�r";�o#̦�2��C���/�ށ�>��P�>��C�u�]�Ĳ"86^4�V]��l�_���"�w��`|����F���X_�6`1p��Z�~�u�t@�w��c�ǘ͇�)��&�p[�	QUKXn�.�;@���4Ģ�$�b�r��R^e�7�L�Ca��p�A�BO8��7�q5��R��]P����us��������������Y䔮	�)���2s���>�~�%��b\�aF]'��"���и�W��΄�;�V�h̴��ӫ�QQ'M+ag=��#m���.�K����0[�ز��[N�{��2��o1��Nͩ~�1��0��&�P�VAm�NI���O5<�9"��ӳ7�()�#�|M��-����8A�@+]L�U\➨��"�^���~�����c��2����&i����&�Z
�-�E��&��8� as&玗���a����:)�Qx�P`�2�8�d���	�;i_�98��p��%:3Ԛ 1�Դ���C���	���
�!������R�T)T�v��%ȴ�LU�p�<��y����8��Wn����0�t�5�Nxx9��A����ؒT�`�o�~�W��n���0��N�n�S.�5��y<w��fM�����!��a������K�SX� ����(�IL�P���r�m� >���!�)B�N[+q���|4�̉�]��(���+��	��~���X��d��%��~�3/�������>���v}&Ӽ���R��U�y#����l�V�t�)-�5��>l��p+AV%����l��T�?��P!��9Na�4�6-I𿠯�j�g'���p9��zma�G��ܸ�p"ve-/��� �/����k{���i�b���E�8�Aj���	�9P#�ݎ�/E�_��d�¸95�����1"�*\���?SC���?��vuJah��5Z&�!c]�)��mfS���ߟ��3oC�D}e�u�Ȋ���C�<
{osY�IK�Cz ��"���q���1�\>0�+�������Ƌdr�Ru�|1�ϐ�3�4��Ǆn��0�'�skȰ���6v�^u�8�(ܣԇ�hs���v��20�Y}i��u�L/
����:���nHx�J�B�sj4H������Ne�>�]^�����'��zGt߾e���_d�ޑ����cMW��i���%A�3'r<9� ���<���r��lr�M>�v�w6w��LҞw$�N��2]~���Q��Eڗ�Y87�B�$g���u��R� �.��$���V�4ae5��;�I�x{Y�5c�xf6bH�J��|q�����"��G�\ʦN�������WY]�Æ
�.�J?�w�&�x�|G�e �nY}�S�R�^�-wHr]a��Z�(��D����"Iw�����J�fO����0Dc^̓���=Ơm.e��v���?I�i�����}�*���H\��Od��?���c��M	J��ͺN��3e�o�פ}T�aha�[�=- ~2)����	S;K��9��@�z\޷�	�k`�'1� Qfƹ�J������|�IcNZ�T�x��2ӷ{��$y�[s���Xd������ m���j�~����W�B=$(����%^)��d��P��ך	%q��K�D�G�� '��zfℯ������W�<�5�Q�s`7�8��F�k�|_LX�
�r�}Ӡ�+Y��p^�a�7u���I>9[�����KI9`�}K3�aQ��Yv���I+�� �U�f��xJ^���F�Xg�[� ��b�A�%�>.mg�G�I;�:up���aM*�Fn�������袸w��|F6�Cs��� �l�(�/Z���M�Z�65f[]מ��Ⱞ֑[�U:�cB�P����Ǟ��''�d�I	� ��i��$�պ��-~�nUG�K2�%�l�Do'6�u�\�]i�__��� l4��Ʀ�e�Z!�����UllЍ�V�e�|%!��1�ҫ�@�k��χL"m�[ZFt)tӬ��tyX��M���" 0�_Q7DR�����E�@'@]�Ȟ���5shj�&���Y�k���n7��h��1*��v���q�-@P
������
bZ8�2I�M��At����|2���J�^ �*�2�|۟/6�A���v6����V��Ԙ�4��3V���������w̡���6����[��J�-HR���XA�L�J�")����~X�1��-U�A�Pߐ2/1SKrc��kY� p���o5)R-r�혅���Gs������R��B}��i_m˻z�+��'2�'�*�7�l��h��=Ԙ�OhQ��R�#q_&�cmP5�s���fl�2s�-Uq���I$'��s�R@S�������=ޞ��,KIPe�B>5[j�i���I��  �x�r�b��W��vR��6�F0?�����x�����{��T�o��5"�j+�&�����N�J3KҾ�*"���jZ��U�.�>�����)��t���K#�-�}�@���xS��`,U�T��g����֖+�2ʿjM��a�ؒ0F�F᡻���Ӓ>2� ��V,�pRa���0�E����-lB��P���F�Q�(�7�O�G����p4;u
�7�V��|tJ$��ˤ���U�C&�
�i����w����~^���C`���M��`Ĥ�`gm��]�n%rd�%��K�&��|bZKƭlA��px�jn�K�9
��ǜ3�Kb���`��Z*+�����k�u��/Q�~	ٽ^��?}��1��Q���y�0j�O��|��ń%�2�����]��]?�я�w����񍤡��/Uuʊ����v��r��S�&􎈽3�
`�E���v"0���ˢ*G:-��ݐ��)�h��	�;Zt�cU!|���Ń�͚��7SY���Ed4�� �D�L3�X�X'l�����%��ܫ���C�&�$��,o0��s/�D��^�ݎ22��ÀN����"鞻���``]�~����߂ư�Zs���D��J1����K�&��3���2�:G9\�+��z߹(]H9�~�B,����԰��j�Oo�N������u�l�7�O��-s��I`.5@��dxeV�#�F~4�F+�}�Q3��W��q�(�n���aBH�-`��nT1����C�G�e[��_��E��W�Q4������vk�g:%����^�/5d�p^̡�rz`�!����ء�Ǘ�Fr��g�_�v3KJb��5;i���<±����2�%��
���ͫTu$�Z�3�.�!~���z ����=`�k��A�g/@�Z���o~��+n�$�L��	7�Ҫ�T5c�HU��ݱ��Ɗ�x��
]���*�>�°�Hq����A��_4h><�@;ۙ����K�孯�pt��i��;��L;Դ&�&�x���n�y�v��Ohz{3FB�a79���?/��-����1�DL����T� ���a�Kz��#U��gݕp��o�����)�.�q�?�F'�l�(�3�ԇ��yr��Y���'�Rq�>�k(<6��=���*�A�lY��*���sǟ{eU��n2e����R�����3�w�7�σm>�n�����-���a�7y�}`�J�j�'L��00�
�$�	�8v��	r5��9���:��M��A *"����:jԷ�9�o]>����H���l��+#C[�4@�15�r ,�[��f}��x�Xܷ㫣G�ύR��
8��ˏ�ά {�ľ��Е;>R�92j);y�nb�㗇��1�Ę�[@�WU��H�צ�9=��)�4�5��O�;9�=�y�aF^���w4��:YYj��1|5a�0l�������L*IE��t��ye�����V�b�.�B[���U�����u ���BFk��88 �Tk|��<����g�gM�2�c˼'a4K��x�ך���G7���v�YY���e����1��PN�����C�%E0;y�$�h�e���P&kM ���c��E�¢׭)�����Zv��a�1P��W�&"B����m����V��	J����\�u/c�
�F�����yO�?��X��%K|�W� ��R� �W�������v���9V\J�һ�eWB��2%Y�J/Ae�0�$s�uG����،��X}�nT�������/\�ɑ���c%���J��dWiE��H�;۴ٰ!l�&�����!��VY��l��vd�ƀ9dmS5�<���N�.-w��Ռ�R���ֲ�B�@`M�ϼ�ś5$ˇ���i)?N���<�D��T&&�mty�R���A �aК�p�$�Q�D�,Y_ +7%=�����~wS�XyĤAe�q��3` NZ�B�!䍽����'8�;� �󱀟��%��h���<�R�)e+#�����U��j�"#
�+�a�u�tl:W�u�ɞ:��2_Xa���o��~T����p�
�}r>S�l�FM��<V��/�<�VN'�q��܇��]���L�WQ� rg؍"�<�%~�ی|{<?�����󻶥�V����&ZJ|��HD��h�'NV�N/��ۖ"X$��>?��L��~�_��d-{*C�N��A���ᢃ�]k�lG�FG_�~��@��D�![w���H��2��C�=�Z�.2�t�uS	�/2���<t7i<I�C�mz��������e���5�o0�����aL]
�L#)�$q�\�K�g�� �U�=%��^F?��QV0d��s��=���6��zf��>����x�<m�j��R��1|q�q��Ʌ��34s}��ve�Xu�KРu&�ޣ-�?by۽خ5�2WX��E��7X{�glt�Q�X��F_%�g��j�m���j!��/�	���i�:}"���ߺ?�B���r�Ru%!RmK�ˏ�������y!� .�����Z�������lJ��Mo��@�.��u���U\@��T�	Bp|��"��>���/ 7kA!�N�C@���v	 *��H���K|{u��/���$��:ͨR$�E&���E���J{��JbW�YtC��?�X�K^}"��x�7���@)�C��M��Y߰g2�ʄJ#�G�sĐ���,t$�N⭕��7�I�I�'�>�y%��+��JN"]Y��D	�x�}�_�4���%%��\Jo�8�J2�MNjN���=��%
������8U�=�r��?� <�Ǩ}K9�L1��Թc��k�|�����S;x�]�q[�|�a`]"l0f�e�\��Y<�h�V��m�j���a�f���IG,RQ*s��N��~w��^�5�>6z�\�a�-/x�Q�E��j>PWQs���᪊{hE�5��U�ck��Y�Ѿ �aO����'u��iK1��Y����{|���Z(P�Q��͕}��It���1"�B��~PK���y��0�+���+ĺmEzW4'�Kv �F7�,���*�;���fN�%��E��3�1:��8�[���OJa�IxJ�*AD���7�Ҋ���8���TL"���������U��&n����M����#L�97���j��pЏ�W�F��h[خW���>D[�
kX#�a�Z#:IU:�C�Uns���n�0��
5v��=B{n��������%�F�q����м�{ +��FG�A��U��ud)kH�Qy�`0�p�$��׭5���?~�Zsg"߸�#n�3��۩�؈V)N��>c�c���m>�jtANr�6 �c90=$���� 4���X�pKV�R��y�&�W����L�喂G��C���)�fU�D7T^ ��s�L���v͟��]>wiE���l�_�f�������K�PCsK_c2����pb��%���`�;�T ٴ�����Hh������{�̍%^��Wc1�X 3�B�7I=��~��qP)���.�Xz\�Vr���mر��o�?�o}`������c�d��a���c6=bq�z\,J�Tdlt�4X�}Tj�h-���Ċ�$vS%���Z��(���%��:l�/c�Wc�}�7�d�	"z$0�R#��S�>?�v��	y嶙�tlSS����h�uR���G�Nm:�~!ukM�>�Sui��t_��&��.%/�����r�i��#�����2�w���*�caN(���<8�t��ˁ�D�f�S����LH��	�$�e�f�|C�w��8���s<c�S-E7�0)Ğ�>�<d�hΑ���d���q�#.P��_ka��?��9�a:{�Nq�m"Ǐ� ��UcLEgP��=)�q:��+硻.I������G}AR�alDh��	7��D��U����{:`���^��s�G�+�*�iU�a���$�德��'�p�f����G�;s��vd;�B�1���Y y�YG�ʟ#*{K)163-�zM�����4
�h0)�,�xV�"sA( G�K�~��`O��]���ؗ�Q��Ͳ�!#�_x��L�۞w�9R���58]�̴�=�Gz�:�\�ݱ���2��rK|W$1w/ N0M�ʴ��t�����t�ċR��:l%������.iX,)��
5��8�j?��̨,�+�9�H���3f�h�����f�W��C's��]kx��hZ���5��m��P�Yu�)���,�{�G�)O�CY��D��~�b�H�T��7��OYP�����;L`��svre۽�p������:`"�+�l>��
�XD�KM�E��\\�!<|�T�b��%0�\���(�`<��O��Y�o���y�:6��N�������S�2� �@�S<�)�]Ŏ^bvM�Z�V���ݝB֥����������R�V���i*��� 
�[�H_�m2T9��86��K<@�Y*"n�iq�(&�+�=�IT&�$b�;ۊC���QbA���,��J*�"f���u��a
g�X~@pb�3<�x�y-���Pg�X�8X�JmMS˥J��G8�R�$~��z�T�������E��(����D{e
䕌x;�8-���.�30+U��"��.Z����E0�`+���x/֚���,nr_9t��E��t	T^��ſ&I�?�g;�+nH�!u��p����W��T��9�oIOl�c�Ě��4�a��6�<Y�14b��H�E�?�`7��CH9�٧�'�Fi ��%������^��*c~ܽiR1 K��Y6��zn8ݪ4x��Ml=�&CF����e������Z����;t�}��95H�.IޤUd�d����C��ka��|~������i�lC��p�V�HΗ��!�?C��6�m�f�(۶�^J��8�`�z T}��B�G��T���8�dm�i��8S1p��Hy����@�2�[�������Àr�U����K��s��?���р�����(�
��z�����Y;�Y�,+V�G�WZ�����Qz>G~KGv׿�B>y��c��b�����ǯ]k���x�!�&P�'�:�J%t��Jb�1:�6g'rb��]�	�.T�۰(N��ban$�O���U˻��r���0؎�v�E��|^��yRs_�� �e"N/��o�3��)�(�Fي�M��z!A�y�d�KI�W�(L��+������J�M��H�Ԡ�s�1v���%\oxɺ?�c��<�J�8�a�L?OB��?�/���w����G�Mf!"����|_/�T�����y����L�I(�=�O���L�b(@l��������_(���e��S""[����C�e�S����f��MJ�}�l��;jKs$X��8Xi=�i0F��%դNh'��
���ɃlB8X��z�%�e�(�=�۪d�T��K�b|lZ 1�'�G�U�����:�28D�T �OV�1�1�:';0o�~d�˒�Z��g����?�%��1��Ylade�U�9t�b�oز8����2ev��2�A��e���6�o���<�ŵ���:{x�"\�$��9�п�rZ�m7�\u	�����5�����څ�VIr�b�`������b��B�N�\��E�vrjt��`?xN�Ơ�e)E���å͊�O�D癿�
:%�
1ꀴ��جK�f�:؍�b���f�|��C�n�X�i*񮹂��I��TZ%?���ݰ�mh�X�Y�F�.��\�"����J��z{�FK����h�5�E��0��IޓA]�"C=��f*���}�*�HW�L�t;͞(�m!�I�5��t�D ��lW�,�0r�ȟ\�ǜڰ<5�j�٥@��_�1`��=v�L��	�����$N8܈q��ܚ/�z������c���/_���dy4����#}%�qF�э�E�����.L�d�bu�Ɯ:��n�q�ަ8RF�]/d͂-w~VES���SL���#t������޵��O��}%&ӆ�{��6�y^I�M�]�D�2?�5������զe���j�M9�z?=��b��6��<��o������V\��rL�1�����k�ğ�8m�Lp���I�[m�~�p�K:�P���`���sdu#��A
�$ހ���j%��M�e��l��U��P��7n�M����R�.v��:�ym����W��B��R��+�V�iik�L�}�x��������s�
S�!򇵇Eӵe�|
�F�U��l���j��G��a�6G���B���E����\j���o���&��B>�.�b@k��H��ڇ�-�P�>��JbW
��=���&gY��d��6�D�}����yacU��q���K�kRN�K����C��7s�U%<���
.&RR����:'=�`��jD�:��{8p���T[�ü�Хɥ�,T����Й�M;�x��|f�ޑ�����;������w��1 ]}Y�V�foX��Px%�7)v?�@�߭$1fgȖ�����@��:���2�.�=�����VQ��F�85Ғ�{��(��tQ�Uru.<z2!��`K�־��G��\Yv4cn�=;M4�I
){�1��6.�����üUW�#��m0#�����ۇ�\�c@I�$	�����}}�����#��}�,���4a��~���w�[]kYJ�4�?��h�a������x�9�d˙X�����)���V �R@V�Xh�?���Ť5��( ��nd(+Z�0�Ny�$1������(���"�|X��)�~U��~�U�4�����rǘ2>��I],XRɾ:+�js�h՘��^yp����2��,M �no�M`����s���a�5*=��F�4,e������d�oj����G��X�ƂR��#�`j0��l�cg�3v?Px{<�!+�vC6�ps���{�5�b[ ���r�8�>r5�^ߘ�	_��_e=S�ݽ�;6�h�:�l$���7�5��?`Tg&XR-V_I�A j)�����Bqch2<���&A4Dj%�M��v,���ȁ��_*������4g
v�Ļ�������.L�}V�JOB�L��SE�.z�UT�]��R��S-��ʖR���Y�D��EwEyZ��*�����iNak�o�C"ϽY��n�[4���.m��V�.���q�chp����m��Vo���J���[�y��Ȳkv����9G�X����7�_�^G_)o�X�M�!�#^�)C�ɳ&���gW��M�5���'/"��D�lY�^�s!�>�\n
��+K�g��J:"�L��9�j�n�h|gS|�*��4^͇L-)E�Dd"��"�l� A�t��s����g��/�*ޤ�[�G����Ӭ��&�G�p�)ᳪk�9(#�~�d�����Â�0�`��8�f��0�h(��G��_W�ŕی�j`qk+�eY���\�#ȗQ��`���"���S�<�{O8�a�#�C+�l�\ �B���6˾�����qS�ܝ�(���4y��@"�#�'�@�>�*��LJc�f�-�l��x��6�O�&���v@KSi����zT��Aٽ7w)N6�8�"��3  E�@�θ��T��zo�?���* ��9���bjj�`%)����'A.]@�G�������q;�M1_���w5NPu }w�Q����;�?�5=^1��ȋ+�<�/#=M_�����ۆ"?�G�i[D$���(@X�8�6�0kl:ӕ�J���/_y��	�Ƃ���^#$�M�k}�r .p�I��t7�?X :Ɗ�.@��+�&�@Ǹ�GJ\mK�-`'��9g�
	o�zV+A�S���zF'seI���b�	a�0�J@�f�����2g�{�^�����L�V)��O$Kf���FJo����d�i�r%(��V �jZ��	(��S��Ya��'������)}K����2�"�Œ�q �e}7�D��� ��w����2/\�F~�P-���b'�JT9�	�s�G����</�	lNe7�pȕ��}����C�)�����V*�0��83BM�[5�`PZ�$0֎	�٬ ��-�?�nW��Ĥ �M�ISw0L7S=Y :��B�v�O+�e����,�L�S��3���.[�z�a�z�l<��������@�bC�Ou�'���븣�ԸC�vW���CGa@i�. �z��������4j��u�[��(�ht;�"��Z���ꦑd�j�������5m�&�xj���X��̰�����8w*�d�V�+
;�6�aҺ�Z'X�Zu�Y9���K����r�"���xs����i��w/���X�T�����Bb��`F�C�L"[_L�����R5gBfŹ )�
�<� �����C:K�:�2s'$lBB�%G/PTU�'CW��2О���"��A��dlG�ؔ'vP] (r�x�Ʋ@�OLs��A���6��<�ņ�ϱOܶG�1z�[H9�<�s�R��M��M_ȿ"p��;9��>�Au��tѩ�q��ڍ�Y���s��?��El��W����~dKK
���f/�m.�m�p��z�)y���%6��)���Yeی�)m�����	��- R��S?���E3A� �h"*w~=��0n~��o���d2�4��"®� kD?L?�昣�G
��d5���~t�ir/�*8W�N��p1�
���nN|�����3�@Q��,^D)������N�@=��ݡכ��Y��0[ �p���W�mz@���%f?�~?K��%k<?WڿY��j�Jc�fL�,�y�NF��ݾ����F���Go�P=v�O��:l9�	�C�W�ɒ`�T0G���A���$�Eh�\3,���(*�Y��$<��d��S���ۗ�h���S�f��T����>���f+��=t ����
$z��!H�o��YQjk��:��ĳE��b]�� ;6�C�i i�����ɏ�M��H��G1�6p�O0�Y49!s�Wӈ�B�. �S?(�wu$�K�p�I��3�`?�h}یK���u|d�������@,D-A�Km�#����\E���uk5���82��D�O�9k�|�Q�)��;4���\s����1�?�D�a�~�������V��٭���9D�a��`�i�?D�1�}�k�&W����▨d/A�;����~�WE@�r�zhw-��E,i�%b����P�x���[��42�tત���KOF�E�j[vaK7`�R�8t��;��`g^��j���y4���{1���4>�j�������Tf�n�ՙ�c��3 �� ٦��~�rjR�HC
��UZ����¡܈3��S�#���	�������:�c�� �#D�E��|��]웲}��H_a*�4�˶�0�A� ���k5��ӝRY��q�u�$���uc���Z`���OwO��!�~���ȁ�-�r���>����͵�
��O��	2��1�(��d��:�����X���o%Ÿ� vM���.��.��H�������{݅YC�3�� ���w�t~)�a_Ӌ&� �0>���G����_��?�۔Wх�(1�������)�{�Cw���>Y��߿�[�:��քgwN-��t��_��>����A�r���M�x���}G��a�n�:K ��o�{����r��7�,���eWͷ��D�#;HC��R�+AW��X��`��t�c�H�6m
|e�C���Ԅ2:"2�p%��*t��,�7\/�L"EQ�P��r�q�ؒ���ے�##���-���C�c�#�b3H��Q�����p�.�U	(���"���ct�Y�>�������Xu'�d?h��s.@�*�	�/�p�����{������=5�l�BĬ{�4����� �Ś����E��c���SKE�0�q�G֠I�n�t.ά���Y�d�s�� ]����b1�@�b����(>w
�7^\O���e0���X��2��	�y�|E��a3]�]��f�塦'��C���|����]4&�~��.����i�����KP
���+���a#V� ����U�Nǭ-p�hy� A�����W�d=_Ŋa"n��aXBq�A��:4l-�߸�����3yR`�$Ga���
\.�����_l3�<�r�%(���N`E�eǵ�zBv��c�<#���W��{=;w��#2��;3��>����C(�C�h��/���^=�:G%���QQ�WJMwƂ�o�p�%<���?A�(����a��o�%1T�]pG��D�c]����idU&.�C6L�����MߦLy �3��d`�I����qeV8Ϟ�і^�֔������+�q�6��m�,�ùR*o#1GZ{G��3��3���GeƓ�cp�phx�e�ؠ�SN���كʝ(�Q�8l��4c�^e:`�Uؼ7����W-�zާ*���7�q��nV����!c�_e�qQ��V�%F�%
�U	��0(�S�Q\�S�^+��'O<?��4p�@���V`��|Ε�㿜����R�����u6�����e�ˮ�
���(X4Yb�d.�4t�6�>��9�v1�5��/{�n���3���(y'Oc��������g(�NցR���x|j
����%}��
"����;�Ft�2z?�[ �߼j=�����|+J-|�J_*�~<���d*�*�1�`�H/�1V����S�7����<#Y�r-�ܟE��!��A<�B�0@�j�/T�`~ v���H"�?:w�`etfO��5� �� �,]�� �?F���	Kw�����)�k=Uz$�]>��h k���kT+E��VК�R
y�Q\􃫣��p�	� >����C�$\:��34�+�������?�2��L�s�D���-�Ί�؃ZWS=��鍍F����A����>���$tU�c�ѐh�!^�Cf� ���p�:u��W���P�"G�	5�հ�(9^�y>Qܘ�gn�:�3�rJrÂ��D���i�b�=�b3j[�������H͆"�9RH�	x�:3t6i�i1��xbH�Z(GUf�jЊebt��K�Iܕ*�?4T�j2���"��LO�,H{���%���O���>�6􊊵,�kr i�{9�M��G�>��!w���UH�t.*#m������Zz�6;-k˓�����a�/��CIH�G��FR�M��vpZ� ���t�P�=9ZӶ�=�����1�;�L�Kxu.��0����e�SD�}Y��'���G��2��G�G�S�����ʊ~FY�NV#�p��,�����e~Q+$;����M��Z[�Ļ�;vC;�r@m�}8O�@� ܀��#�1�dMJ;^����qoR��zG}�x�G�'�0k>��EQ���P%��@��bkf�~ŉT���v���'�Bڥ:r�̳��B�^���@�SG�O8E"����cι�aIN/��ȥ���44���)
դ�k�pf�U��������+v��8PI�yGga�N2�C8�a�~��1b.˘�)X��������{���K��ʑS��|
a���x�t<r#��zݵ)m�XL�tWzЈ�S�%!�,�ȯ��<>��̢���f��9ꊓ�D�_��=5�x��y�<�k�戮BZ�T�:W���$u�q���^%��%�N��ܻ�]��@M��I�S21rK<
����]��{�?���#$y�1X�7�]��z��,�9��&�
*�TS=S/�B���gx����q��3�̧��g�dt�������N����E���6�(��^O�b=�#�2[����掠�e��-b��9�?o���_1�y$�A��$��s���	4���b:��d�X)��5����^D�%�MN�t䟛���i�=d����:-���C���[t��e�ym<���f���&R3��*��N_�?�i���#a�O�x6�KE��;q7�'��݆�pzI�"��ݣO�C?�ˈ�[ϔ ͞���yO W�G=� &�T	�No�;8�z�u�FI��� �vaBT�HJ��O���s�W�l�c�[ު��0��y�jp�k�;��S��?�@�t�xBwCt����0�z�� 9>��=w�b����O(ex��!J�����*�%�A=��l���:D�.�2}i���-�P?@:�[A�0�.�a��!H�s�!��;�d{�a�A@2�f�����J�\/��A�\�R1�s�c�������-�!�G�Y �W�t�X� �H��r�iyZ`���xS2��i�4O��oT�L4�Ɍ*��;@t��D0P��F�d�E���x����Q����g:��{�X�bc7&@w��·���������J,L�� ��!z�Px}�a@���y�==��Sk}�I
����� ��t�!�U���������U�$�I%x��5��5YeC\@�V6�K;�B�,��Z �x$�H$��n�/�"�	oi��S���r?�����C�?$�nd�n6��8��;�o6�K4A�fУJ���]s�/����?��]��-a:9#E��#���Q�����d%J�.V�K�;��>\��"6'ZrW�+),��@jJ�rC���D_�1[
�nޘL�Sq�}҉�6�B�]��H#�ca���zVh`<�(�X`3*�ef�Ζ�~Ag[���^"�ax>��e�"��P�8����`w%8W�� OS�Ƭ�����-�em�n�^�*L��k$�#�?���}]Q��fF�J$	�?F���z~=}�V\��(�@RV�u`@*�C�w#~"�(��|f���~[^�^]�.���p]��!'�B�8C��_F���ʊ��l�;�rqŦ��7h�U;�j��4���C���O�'D��$Lh��ʆ�Y��G��:f�;c���]68׍�]�!��o�8�B�k3��W����+�6S��6M�6N�t��V�� e�d;��Ӓ��N��3SZ�L��95c^�z�H��y�0��R���_��1$O�KpU(�B<�*��hlPnP�(f��R����/�V爌mG���ǉ$����%��Βb(��R��v��>�#�U	cm�|�T�S�4���xO��HD'��]�cQv��l�M�x�ʘ���
i\m�z�R�����m�2ϒڅ0��'�x�ؽ���W�d�1I���?5��/�d2�C��($SF2^�ty��S�t����[�8�{��#�tj*�KB���,q�+_lA0��`(˷ah�<�si2BH����*5YE�`�f�X�x����Z�V:ﯭ�s��ֶ⮪t8w81=��<s{KPB9����U��o��  !�eA��1lf�ޭ_d�ﾁ3jw%�J��FMFL��_���X�
��s@�I�/�I�"�&[A2����r���a���-����e����b�{:��s�F��K�\�Ʃ~9���ed���78N#�9*>�u
ɭ#=�nb��rpr�����n�k7gD��KR�JXM���k�����}�/Y;�U�(f
���酄�-��8(��pwwq-(�H�y��ZΑ+��3V{J.s�gOvN���_�{+|�<��\��c�0��r_Գ�^2I-�P�$�ap�k�s �Л��[.R��K��4q,t�藼��̿Dǹ�/����%1���yBV��yIN���
��r������%7�<cS���ŋ[~A��52�f𵔎K�m9�[��n>1X��l��XK˚�f����II#|�al��t����8�m�?�,����`� (34���xy��dgv
��O�Ԇ�{�� �3�#�Q��/��{��6���o���&HR��������}�T���x �,�3�d� /�s���'����G��q,�O(�iMA�`H�.B����.9��GK��u�Ǉ7öcf�GK�Rv�qn�Zo�6�Цz ���ˌ��~�{2�ͻ9V�~2�X�ۦ�1{�ep���bo*.��XN$���x�(�?��ʺ�^BC5�۠����+�A�N�m?��}�Qګ�j�<%9�V�*49����SUF[&ҡ����./l-��9Wɦ1�)e�4���Z�M�bcƻ�x�t��.~�D���_�n{3>{yn���1t��$0�+}�3i��_ǫ0(����0��!E�cru�95$�U-N&{�s�H1��"���\�T��n�&L%Z�tk9�`�-Yݸ��/m05�>��]!3�x��m�q��&���g���h��Uy��2g�@�K�DE�r�͝�Z�-�1B=��?�!MqG��������fDi	�ڍ�3�S��Ft;�Q;�Y��8��#��R�����?������8#$���
�'�{
	�0�^6}I�>�}�e�z��.��@��5�j�:��-m�_~:�09&��L��
a�DA,5\�b�\�_�|�B�>�GZ�Z�ov��l����B�{�<u��%w��c��y��}���l�3J7�G+��;Q	D����0x	��Q}1��S�H��9�/�dRۢ��^����(p�i7 ���2!�̚���MJS"�r�P���{>V������U���a춂x��Nw����D��L��xߢR�f[Y�f�g�~qE�Ď����qR�xL�+�l$�M��\���ŭ��Z4~���w����N�w����
3(Jyk�q:aG���$v��mǄ�K>'M�MU�2�.�Ub�I�l^�Z�͸�XP��Q�e�D+�ҕM5��p�f'}߬�BU�9��z�S��D�������lGw��*�J����^�EL�{�z띳���"���B)ou�dV���) �?�,�>}�C;@�XiA�c�o�Q;}�W�<�>�3z�op[�g^=�u�6X�eX%` �	vC�fI��=�Ǒ�.XQ�k!)(���.�M~V��;I>�o����U����l]یV��S����F�
^Z��r5��2��.\���zY��s��D�;���OqѨ@#R�AyA���M�A��QI�KJ���0�	?���P�U�5��!wɡ�{S�o���"�g�B+�z��=0��8��J�Mo�ɀ���a�,�+Y�����W��8��*�b��LO�b�x"jo�^���z6��I3�b@�L}�~�������g0!�ӥ=Q%���W�I��{V#��o՞8����lvv	z2�F�JA_2\��<��{�Z�Z���=��<����n�R%�\�Dĵ���`fQ桜Cyg	vLO�:U�p�&�^9�h�my�.�e�+���׊Š/�@ZD��,R� �<ĸn�.�RP����/ �fm�5��!�h��Ԛ��W���΅��_Ny][���w~�|�ŃL�R��x&e)�I��Xi����|��a�|[�=��F��X̅���������yIPdmv�����&�ӄ��%�Uϥ�/-��&�m~*�uN�Ļ��T���Y�0�̚�+���Ч��7�v|��H�W��L2@��xN�?G��bȽ��FP�����4��L�v��s���z�
�e����wR�A�U���K�������L(ݴ����(����	3���˙�A?*`u�a�y�)=�%
�`���	ꥺR�v�Nv���^���=h�`XS`d1��^���-�s�'H��?4JDAk�rr¬�\?<�B鯰�઼I5����t���Hl��Ue{@�Z�!6�"������wT�{V�M�<M�L�,'lQ�]�'{�y��~ϕ�m�/�����d(�c��!R  �?����1Q��N�!�aI�>����~�OIW%�UyǄ�o���K�\�-�%|ܞ�1�+=�~�Oj`$�U�U!�$�]W�mQ��O Ưj�jĬ�=���V�>��XT�H�74[�����~���v�.�j@4B}�V����)����E�";��(��c`. 1�Z�,ɐ.=7���s^�8�;ws�����S73�&P̓GR��,$�9�b�;7���q��~��`'����Z� oo }�*���n��vF(��tL�~ '�V̙Ĵ��m����i��D�y=�xCI@��%S˼��v�E�s�,Y�fq���	at!�'(�eA��w���1�c��\ha�NI'x���n����}x�[��!+6�3�4��uk�H�DHp�x�X�O�k�w�+|@ԓ+J��_�~�",��P�:��,��~�0s��	-6�ߥ���3�s�gv��O2��-�-U'p��B(�Cy��?`;H�>vO詃�����l3.������ T�c��P������T�������S�	�N�A���1`9l�$+���k��Ge�����MNr�a,���X�F]ڄ�		�@��ݽ�L��2�;?�l͆�7�k~�@���>"K�bNO x7
����M��#@���O!��|�XQp��'�0?G�d
W�Tw�i��7�J�����J8�[�/�[d����o�� D@�9�]���c�H�?�c�8"�x-)�o�G[μ����7hdF[oGC9:q"�"�����e����1_H66�l)���#��Ď��ޔ^�s�g*���
	�k\�u ��er���`�e��B;�"�I�)c�ܚ���9i.j`W�@���xF����6cP�]�'��f��e �+��&�V�c�2/����F>��_�_��d�ə=Xx���`|\��f��A����q�?	�f����k>�q���r!���nh���:����6�n�e�!�N�/�'�L�C��˭�1Ȼ}����Suq�t� 㷮$ꌠHe��|u:��MC0�/�����C�"?�W�IݥVB�|]�v��>SPr�TnQ7OpY�ERx�eۘ!�{ �ݯ_PT��Nre~���2��7�9z����%�\�)�I��l�F|���m�[1(�yz؍
-�����T�]�}ڛ�A3�#����^)�^,�����L�}�i{��P����U�- I);���F�\(�C �����uh��Kx^��9��A���5�n�#��)7}ٓ��&J��w}wU�Z����]"W[u`]��(\���G��h��t^{�24��!��w�ȇ���-�����I�-"C�@�p��Sʁſ+hdD�{��Kn�5xT"��@��m{O����q�>�	r��j�@�} Ó(6+K[W�+�]c�;����l�I���,�&Lz;Z P��ۉ����=�r6t��(���tή�vʟH(�j9�L�Ϙ�@����[�����zf
��N����F�5!���#g�I�aJ6���N.kM�����r��HQ-�͘5_��Nc@�ۊW]�I�M�ښz�����4�G�iM��I�ގ�ex-h�T��m@i�e����z��ts~[�WJP�C����L���P�͆�^cA�G�}����ò�ҩU����{G�[�Ey��1�Hg�J�BA�e%��e�%0x0w揅���K�}GƷŬ_ċt� ´���r����!�B�U%}�cׯU_`/b�K%+�b�>�C#��*˯O�*6Z��[�I�ٻD`���Z��YƜiƍ�B,	�a�'�����2dF5�����l\zLplX
0o+���E�%(3~�ߘR��$��W��̓�蠑ֱr@�e-�4���������֚0v�-PS�y8D��
U�Ⱥоh=wN�X�v$95&%2���[x�{��L2m~��yQe�!�n�N�=H�T�E|�G����D��ǝi(��Xm�0l���k��)(�b$��.�_�6.�G�����|)���YU���8	s�)ē��W��x�	��>0���bߪ���&�<�O�ƒ�m��Ύz��l:�t��{h,���47����Ӆ���3D4�w.~�џt��̲��-���W�a).��x��I�;J���R�њ��B�<�ɞ��Ξ�L6n��.G^ʴ�~P����$8���Ea��v�*u��Ji?F���1yi'��l�p���S��a���]ɵ����水�6G�Lڑ>�=�������VY��ѯ��#&E��c�5������?.
�Hw�݇�OӀ&!<	e�\��2S|R�
猯-yݛ����׵�4{�וtj��o�D �7ʰ�����<<�RF.�K��%ȥ��-(�y_�+���$,�m̊�gp�
\�8N�K��Ev_mvq`�8�M���4��V<i���۶c���7E��Yq���nSv%��vm���.giJG�������$"�E�u����ZY��,W�t�G�ב��=%k��w�\⋊9;�4�e��;q�0��b]�F�a�!���k���z=����םۯ�؂r�a.��`ZP���H���Ӂ�����β��ߤ��W���=�e, ��0�5Gy�j跤�(�X����Zz�����	.�X�����w�D�tP~�I, ��/�sG�ٷ����,�)N���lL�n'^�Wڷ����A�Qh�i�q�>h$+��\���&/٠&���#J���!�>u:ʂh��T��m��^�ϦXw�5VjH���a�*��5�a��	0e���k��}.���t���}$Hٷ���ӽ�0�]�Q���r6�<g����5'�2_��b����H���GZ��h+��g�zF��h�i	%Ԯc��fC��uǦtBް�,j���P���I3jue���u�|�oz;LM}V4��ud�;2X)�1@N<�������V�v
 ��ݿ�����0�p�,F;�M�5l�<��3�R� v��w�R���47�l�7m��Ĕ�i'�l��]�$?W�Yǂ�}q�þy
��
�`����&^d�;6�l���6\�dÖ�Z4B�NӠj�k���M!��(4��4�{�(�M�8��l��F�R�#�/�����
2�bL�i��=M���1�x����i���
�\���TH�	u��&��29AͯAe֭�1�*	���9�B�<8\
�]��":��7��z0g	>���L]�w,�U��:���^1����}��Sa��ew���zor1�;J��<?�ۺ��Py)y<�����o�����M�NA��G�9��
-�F�_u��8lR������I;�-�p�S�w�$̄�>�4i]JHH��]�D[TIw�����CF4k���`��1l�Ĉ+�<��V�M��֐w
@�2�ۦѝ�Q@��U�Br��wa��g�`��D4�d��l�tן� ��D�'��P��!H�hܲBb@�h�W�@2wY��c�\O��t�v1���n��8�B;�;��s�}f����&O������v׵��꼚�5�v������ɞ�%~#?3�(�.1��wW��e�Lm��b���4�w�Ke}1����R6����m��� ��*�c�P�~�|���!��rM���(2�&���XX@~��GwV�fR�HU��(b?l����[��t@X�l��ȥ6�r�I9d�>ͬ�&ڠ�zМ�X�'�Ms��M��ow��	���ٳ��k��~3J�BQ6ڣ�(R�r�� JQLp(qf=�I�7Z���=�nqr�����c�~r&Rj@�e����c�P���Qg��)��l�xއ���˃���� TC�+�덤��o�'SV=l��\v���9��:7ǋ��KO+�9�/��yN��q$Dk��FP�}Ξ�cfrU�"/ [����(ԱdB7�-�#��&s}"������F�9��/�R��z��7�������H�-�
� ��<8�{*���W�u���>���u8�J%<�k�\��@��x��>��#���
�8 ����O��/O��dVDiMi���q�<  ]j}l\����N�u��a�+� [�Y����H�rEc��䤦�L ��B���'��v��
U���� �M�&>�R)(^yж�pT2<�o�Ypf���4���dZ�@�[{�|���5sغ�d��T��#�(���K%!�Z/>� ]� ���BTNPqM��u�_��\9�������K�$�� x�(c,1�6zӡV�����9h�Mi���'5�����b���4��Ivǋ���Ϙ	 ��y�c\oi�~�$ʡ��L�����ڠ�[�n��&I�l::�����BWq#]X{���P*�=� ��5�!�`D�u�7�����7��u"��u�F��=�G��.g�L��;�,���[J���4+V${t���-�Jd�%mN���
""�A�I:G��2V\�;�h�BÅBǲ�f��L�R���	|��׬.y�1����3Ƿ�E�i�Y����S4�n[��y5»�N����v�Yኑ�E�82iE*,u�߱x�3�=��
��-ץ]v���ᡤZc�@Zo�>��(
���ҔN��vSo󈟂�F4p����zMVb��ٷ"��Y��P�f�+K�%�\ꋘj.��{J��_�i�^<���8%-r2���������7�4fYr!b��:dn%+SNT&��b�4 ȑ�A�![�zէM`�_<�▵5b�����K\O\�����ў�/'����of�k�0�/{Q�r̗�o�R�3X{��>��:O��phC�+�7��~��s��T���7�1�p:�����@	�h�挨�u�U9֣�q&�Á�y��s�#�ޣc���)T�e���Do�|M��r��4+A�*(EW��8Z�� j�0x5I �����;���052��.;iDh<�Z�~���WB�>Q һ@�R��2�8�\�����`��G9L����7n#���.���9����#��N�I�QJ�g�ol��	�rw�3�hBwu���ߵye��J���(����@���ïEU�����7[���v!2B��N ^}�Y�����J���y::�.�o_St�R{|:1S;Q�横��
`ՈW3 ��A1���X
:9��3L��8�,��npV0b��@� �7���[�7]�Z �ؽ`�Ի/u��o�# fe�i-�
ƃ��4��'kՀp)�Eu.�eE�K�[�*>�L+\pe7�h��V��p '�~�x�0Ht!�Z�(��
�m�#z�᫩�`#�6*��{��~��9#S|�FY�/%q~�t����u�C�x�H�?sg�1;
V�|u�"ˢ��1��f�̉`�~�e��;�N<���.D~R�\d][#{�Z&����J-d�Gϣ%�#�_e4�ޞ��|�0�L"�0"DGY��&}�� y"�_ʪ�ȴ�F��7P��{3����t�x�M��C��2~�� Ki�	��r����h�vL�S��p�
N����۷�h_��Ox
Е3|?��b���XT� ���:��3@�|^�7-)#�E!��l���ȁ����]� ��J�ц�L{J2��j�jw\NL��'�b�V4���}|��;�_;Y��D���z��FH�3Թu6���:��pɞ�hB���b�a��w�G�֍�|��#��`luޕ�[�RBI�q��k�=G�JE�tP�k��`�Mxg���c��:����M�d�?%���FR8��=�{f��'5�鶖��<'U���� ���2tDz�	r �<�eP��:�'��y&ѫ��3O�����ו}9\�.��eV9/s��G^_=��%���/<�dl/�=�	T9]�Ov�(�^q�2������m8ps �{F� N�Y�gz�%ח�5�,����Z�>e��:n�]��bA����.�E}�x�W���߾�u���.��2�iE��&X_�VP����$ ȜJb'z'I�-0���io	/�x���>,,,�Ah#c�{��m�5ʵ���Rf�� �vw���V|Q����υ��$�TF��v��0줟z`��M:et�I��aR
ft��qь?�`Ze�ж��7B�;��I'���,�2�4�Yf��2��*=n?�H��Hj��}��J�{���]@����N�&�G�S朳_�Gk����5�H^l!硹9�v�͞6&�w	v�|�z7�މ))���h�aԼA�z�h�_'H�:W�m<�Y�/
�}X���H�?�Ōdj�iD���=�����qP��E�M��_�ǜeG�s��h�H�"�;[:R�����ň�?��QH=��G����}��)�K&����N�;��U5�O�0RSK.����!���j��*n8�|�ͤ�pAp�#D�3>��%��Z�1��J�3)�M��yPIW�F���z/읗ы�x�ZY��
G��!�� �-�?!�} H��a��C���m���k5UPϤ]>��N"���Ƚ����$'�̣�GbRg8��g9N.��lR�ǳ �i}�U�_�,Z�G�����<�ն �c�C~/4l�הe�o�Q�߅dO�C6�S#������@�>q&7���}<BDҎQ�����f����}�9����&�R�
O�"�#�m�6����c#3��_}ML4����})�S*ӻ�y:h9��<��3d�FLr_~�h V��뭐x&2�0�.�������Q{�NEj���Цu��(�+��H�6����+&2�46ǝ��5@G�=�\H�|��P����G0$$��ތ�c�Y4� ��6�lpې&�u���8�rz_Vc���m�:y�IB3��'����y7c��-��N�)r�+�V��,M�B��fic���\���hC8G���f��V0Z�<� fAGے��L��[Z��JD`x*���`���N;!y��>}�Ћ�e����9��;��T'zz��%r�j)X"�T^Ƥ�ś���f��C�gvfsPק�#G6�q�C"tce��9��^Eݾ����2Z�����q���:�/T�2Rw]ֵ�`�ܥ�xO6v"��NLbC������o'��]C\'���M[UN�o�<�@��n�x�c�8�xn��&h�+|;�r&����`���aź��sb�naX�t�o~��'�����VS��c��7`�5M�Ŗa8w̵	nX�`�Tf�Pԇ%�nn�5�W�ՠVf�Xx���}R��w]7�N�>K�Uq��¢�g؇պ%J�̏����|V�mF3� ph*p���$�qG2������m�Ff_�-A�ݺS37����Z~H�c�x��?�D�L��;�c֭�c�^�8��g/�x�au�ߺj"Gu��3�#:�̧��҉���c�##.B�Ȏб T��_��OTZ�̷�O���}�^Y�U�z�^È��n����}giM1�����f���kn��C��1��3b(u@c c�M�`�����]�&�t�R�$��`l���:1k��^
g�~���Q#l�+�2ʑ�cQ�x�Sf��I
5�,�g	mCrѫ�0�0��#]�OZ$��@���TP�����9[�Bb��Y�*�(@hV��_`�~r�o@����](���n3��Gu�,�q<��Ǚ���l!M�<��[n�� )�O6����.%�3OjL�¢��۟
�%b�.7���`�?mNL����Iw4�����v=��՛s&�q��ע��'zg��Ɗ�4����ʊ�2ǤY�YP����X���\�tet�$7�'�ȓ,TA�'An࿻�*�g��ھ�b���-���r���M�qG�7�j�Ը7~{	�ҊR��7v�>��Yo}��\�� ;��B�T�EEҳz�p}��@�X�X'!�k�j�@�T���R)�Uq���f��V;�����K�X�]��k;G��sl��������y���%e��bG�@ �nVZG�f;��fhp�9X��2�)��8&�!������T�?UL�[4_���"�w��8{�ʈ�����E����G���0��o�/�co"���qTd�7s��������BP�O�Ӱz%c�ڶO�x��H它�q�֝���H�B�*�'3�����I��1OJ���_Nrp�ᾝ��ڏ�Wo�V*����$�!Y�l�����Ѐ_�����(�R9d@`j8�� =.}|���x;A��p]�b�vt�ٗW<��A �����鯤z�;&!�E��%ayZ�&w�@͇�����]~�Dl�V�?���%}pZ�#ͽ�q~�аD�u����X�Y��"1e�XP��M�QC.��dI�~*x#s_l�C�&����	9�ܷ�P�5���{/��#�nl��K�<��!�4��2.�r^���kkq��?Viߐ��pV�D�v	,��mY�V����>���S���V�/��#4��Ez�����["�[���k�Km�����h����p���nf���
_�M�s����/���3Ŧ��`x_������,l���8q��+����c�39&�?���s��G�gۢ^������Z��z_L�Ti�AtA������ts�;z<V��k�)�m�S���Ӝ�W,�F�I�v58�>�{�S��1s�"<9NQ�zj^~�7�܇U��g�,y1f{�����W��RC�sO6o�4)����}#��7�����&`�m���B�~�{yW�'�l4�&?� �j6�ر͊�V��!����L9��+���B�!�l0�Ô�m����F�ZM'a�������5!�'f��h��껈�_�����c>E�CP���PF�m��(� �М�����^�j�X��E��1�>�߰�a�P�2��~��|����TսB�1g�K�����Җ�r�/�#|�~
Y�K�&7��_��S�S^�kW�y�d��*��r�<��/.UA�oFV�����O�z1����T��H�|��ƌ�Ih Ɩ��d�N�9z�J�2�_Ay�`K��w�}����'�_2O��p5���;p
��9�PA@���9����s"2?�[�,�;�}X��d��3��� �)KU�r�<L�$m����י�#3��� ��:�he�j�.��JM�0��řP3�>ē�='wY���5#�
R?E3^".N�{X.�A9��ә�c
!:�O��D̎���F41���-�_��0+>X:��q1��v���X��Dy����k��o}>]lK�J���>��v$̷Db�1���q@u��R�vo�i��K=���	�� :�aLT���:_<�M 87b?H�_��O@����(�k�&t�>,�:=��l �G�g#��n��_F_ߞ"�A�߉����C�Y�6�� �������1��� ��}]�I�'����h����������V0Ұ}���9^[����� '��r �\a�{���[���?E�<���-.�GW�F�C9��nvk�I�����qOT�_��u�yא�vg�D�`�w�Jk�^r�=Q ƹf �(�^�0>V�ؽ�� q S�N�W�>��Í���Fֻzina�;���h�^tl��+���$+���7W&*Jk�R���T��-�U������G�d]��R�µ�g�P������n{��C�9�=IISN9�Lq�Ӑmj1��͛�?.��D"�z�#L?���R(��(�~�Щ1`J�T}8��*,�Ӂ+ܜ�i�5����C}���Ej�	�Ց���v���s��ˡ.M�䪨�Y&��="P+�ӕ6�^*"�ڽ.�����

�UQ,c�Ѯ>�������g@�s��y$���l�k�bIWA3��`�R鑲E�/&�V\�`!e��\�[�J�Nh8���-��T��@��ʛu��|fIm��Mgl���}��>�Pg'嚕!�>�7D�y�M�!����r�I�Bq�I��^������X��:��aX��X]���xÝg�	{f]G"&�(�%ykɑb�)���ˉ�^���Q[ȅuW<��K�U�����q`:n3�n��h���A���F+�+���Y��qMw��c)Ņg���mz���zЛzވe�a���8V>�6}���K��Ʀڥ�w�we�t�V�J{;�c��z`o��K��Ќ2)�]I�*H҅������؆	���˼Α.l�E!��EEʉcn (�L����y4�q;f% ^~>�a���t|"�dZf���^�U��&l��h[��d���]�9��vF$��"�𙖻r ��p�<�H-*�S�`-�,�Zds'���JH�$5KR�߅-��j�K9���U+P��='X�w����#���-w '�q	7����I�!I�j�&��k�p�.�����B�^9�f��H{N�uI)Z���Nh�L��ڛ#Ѩ���:�JJmU�e��ݸ��ƥ���7����tLyV�����F�)^��/�����[�߆�����O�i������+���]G��5Z�@w>t����� �Wʾ!qjQY��#c͋xF���QR����Y��Bd��T����6fd}2a_�|lL���*He,&�#J�����|*ӗwh/^�\)�S5Ы:,x�L�8�R)�.�=��cH����<]p}0�dl�|;�U��X�0y{%�2*��^�O�G�&h�!�2ze{��:�\f����[�ӻ�q�����6H�˲�K^*�ɉ�#i+�1+�?��H���q�x���σ�k�zz�8��SqPX��P�5���DR9վ�ڊ�cꡲ\R�Aܖ�Nό���쟐����R@��wW\C=Η#��?'�%�<׈��ۯCШڛ��Xiv'D��8�_[��(�iF�*|;Ѵ���~�+Q:��c3F�PS5;�3��D���r}�����x����=;�`)ǔ�vY�ѡe#��4*,�[͉���X�^43�/Y`��lA����˵�d���y�gk��&Yo���$Ґ�9����J��z���8�{�g��Q�۩�2K�D�����b�Ԕ=gE|�Tݸ��x;k�f�3O�6�W|�[���:=v�Ub�P��էB�>��o�{�Ğ+q��00��W�:x@�L���������\@�9&�nt#�����t`�i����^f�Fvu� �q�7��d���d�)5�>�U=\���\�_C�\�#�ܦ��?�v��K
���d{��@���E����$�
�J_�"1��+�%�#�s U�3���j��������X���������oR�k�xʔ��z6�Y��r�Ǚ7�77Jh��jݒR�^C3ҷiD�d�����k7�O������#R�crd[>p��6��ð5%�|QS<����o['��7�(�=	<c�5�kZV�F�_�Ѵ��A�uY���WSm�Ѫ�2~9�͋S>���1z]�93,`��&��q�V+>/��=��gD>�h����O�Q��DM�P��{,�5�Ͽ���}�Π�,�R�S�j�T@@J��5 ��ô);���_/�[&x�	$8���tNZ���$"!��8�Z��[M��"���*uyxU�{ǆ&gJ�����2c���4�>���^��0	r5��;�sh+�I82F͢N\��~;�wX�� ��_��T;ۖ_��w�HkweG�G?2���o%��pX�w����5����^#o�,�� <Åɺ�ԭb�����i.$^���7Bm	�h��%Z펣l],i5	��8<�#�gȋ�v�Rj^
�}G!���l��?6��T15���zj�
��p� � ��GE�g>W�z)G�=	�3	3�w!�����@;~:W�� �7���A��*
x9Geܷ���W����������E�Iݞ��ꜙ`Vb'�[��NJ��K�ǀ���ӜLSO�
�L.ҪR~����APVwm���)������mh���ky��Q����\����uZ��n�L�O��d�Yq�z��Zjs�R�(�؇Z�7ی�xw�}~X��� �|��𼉠Jy������<�S�<�F�5)�h��錢��?�s@���y_����[e30�#;�8��'T�"t��5�J�]~�~}~��=�$bU
��CW �	S!�?��H*��*�e�ت�D߫A�!��}Ɔ"���@�\n<)��0��7���\��Q5����e:���>l�-��Zv)��U���ؓr���A@�~�184�����C��^��øQ3��o  cIB�S�96�,Ҕz��Bk`��LЙXV~��������muT0��������䁆�k�p�p7�#T�����C���u�خ��**��q�`��(^�����Pc	f��	�%K��꫅~/8����u�nO߬,��5�>4�mI�����)+p ;�E0V6�~��7�ul��Q��}a����VO��!?�1J�W^�|��D�P?M>DO��BzR�}�EK��=F��%���bm+�N���Өp7��[�=%���A�Bҡ������~L��g \,�b*b~E�ֻ�p�A������SԖ�#�)���3e�Tj�m�dn ��d+M��(-qp�p%h���o�cW�!�b�0�%���~��ϕ����	�B|����`�tã`�Bk-n�s��� w�q��+;��5���G[O���G�R*B�n@� `��"T�������c�E�i����M��)�k�(�f�ΟI*`��G��-�v5��MG�4^����D����� �6N`Fh�� ���қ����7{���;a���[=�����d���	r�6M!�(���v����G�K֠�3QQ-���B���k�	��r�a.�6��*��G���E��I�y�?��>_r�n��' w���o�%����
���M����=7h�b|π��k�7iBYe��W4���2	�>�wUa�0�
��WNXڊ,t���=�b	�
�h�|oڌ 7D�۩�mGN�����{��Au�
��Ȩz���PV�g`��BJ�������dE��N��L��
���ZZTs������eA���52KX��񅽣`=���E���5��wl$+
�����cM�GU+���L�A�r ��v��h��{�2�
ra��R��d4�)�k!1��hY���؈8��K�<�=0�dZJA<�0J�r�ʩ�[ۡ
~��_�O�t�[&�E��B�<e�L(�H$�\�(O|W8���.�ݮK|���&ze�3Q��*m7�  �\Yl����ڳET�$��D�K��qU��ַ��*;��h�z���%�"��H2,�gt5v�8P�i����&q�J�6����Ȱ��H�jW����n8N���힐�����OUq���B����_Mf}+�XW�
\�+��w�dy(�F�`[�%@T��s�O]7��x&�o���@�[���Zߩ�+��5U �+^x�~�&)x���{PI�ܢq�mAR2���D�>�4>;H"q���I;��5n"�:�G<�N��Wh9��D�U��Q>��[�e����-���OMX"�z�.p���j��ߛ�� �E
+�f��� ��z��C�A�p�����oi�/���BxvW�Ї����w�Lv��7xW�V��t�3�%��eΦK��t10�餽>�OJ��������y3̤^�y��Br��5�W��e��6�`J��+�{S3�<��@f���L4n͘^\5.8R�#J�l|�,u0_�QI3`�'�Yr&�Y�,����YBpr��W:�v�u�>�6��/�y��[�b���_+��Y�A�Ӵ1�~��8�$}GHM������@������v���H�V�H�)��+���7{�N#��;�&@�}��y�)�y�{�up����|���{��	�����ԩ kF�g��3 �	��W�
m�?L'��h���:��c���4L�F7Z�	q6V�tY�=3O����t��zP�g��������M ��`ć�ǳ���>��ԝ��M�.�^�>����&,�2��5��v��g)����g�t��>1�"6S^��˃(/^ȫRUv���L�RT i�FВ)Ǆ����ۂP�
�x���?����ۯ����v9[z]�b��D���R��0�s�YT�G6GB�I�Z�o�yR�G.r8'�j=:�ogRx:g�4�O*ՉP�����y�����K䐿��f�(;(N>�(�P��Ϧ頠R�աf��oW52m��*[�Adw'�نb/�[u���n�5g�"t6Iv-�x���c���P���B�;չf���I���ߏ9��a`��o�L�Θt:~מ��Ȋ�	�-WU�]�.�ށ�:�!� �_@�|��'}v\��Qk&E%m~��s����bH8w����bSF�`
���!���okj�TV�GfNd���$_C,�ZXk ��O��!�d�Z��g�1t\��<r]롪��]Y�oq|�:�8r-a'Z[�0�H{�����h� 7���j����;Զ����{(��(ib�Ec�M���{�T�ǭ�1а��H����6��o� %��&���4�*�n�]�3,2{߅͑x5�M�?mL����0�#���� x�S�/��W.��͐�;��b�ԙ3;q���~�h�?=R��͋��	�x~�9����mbf��&/��;��m+9O��Ȳ�w������W������
�0��|���� 	����ho��C�:+�Dw�^-�u=�8�������w�G��m�� i�� �DU��	�I� Q}��]�{p�m}ki�32F�r�4nG<"�t�;�M(oڋ���-=0]�v�tX������6�A4��kk￧ɵ9w0�T>�+���!�B5�ގ6H:�l�vQV��M/�&D:-��}����l_�m��<$��	L�p�Ts�ǯ�Η������=o�2N{��&�a�Βt@a���������Io�~��\n)y8��DXʘS�&�6J��ً���"W�����ȍ��ҥEV`*���-6�}�b��E:b�Yo���}�s#�L��ځ��B����4��8�˾�҄+���o���u��X�K��6�}�^&�%{���� �\Z+\F'Z����s���k��Z����y�}���6˩;����~��K��ŉa�75����1�eJ�kC�u_�z1	[ym)�"�I	=d��s�*$�^$t��u]�D����v�&��(�Q=��b��fT]!-(���Kͬќ��̏y���y!��Ki�1���e҈	�?�>H?}Ou�T� dn�5&p!�#[v)���vw?��.m!�}�n�D��䞭)#����!�)ܰ���M�1�����4���I/�:�&5`R��t�͇���P�7��%�Fy8V%�0k{����E�Y4/��໠�A�vG��jO�V�5$�}Ak\y���?����,��b5*�xɒ��~j�қ"�s�_@2��+�w=��%�L����*S�>&
 z0= �|��`�#���ߩ���c���>��ͮ�E��0$H�o�P贉@E��� ���~���B@����̎�Ӿ�����PC/-u��:�o��q���{�����k��j�Ʃ-�|�j:�4��J�\k��ܘ�q!!u�|-Y�4y��]� f���_.���\X����xU]�z�ķ?~̣	D!2�b��^I+��&K^�;Er`��d�=��E	��~��sS=h���DK&L�l�� R���:"�|��^wpl�}�Y�fS4��ߺ?���Nl�r�C2dHk�?gCE[16�6��䮛N���9t)|����@`�\��ڼ�BǾ�\��/mJ���t��]ո�5�_��F���u��d#�A@�	\FPK�:�I�=��ˢ�].��Q�?ܮ�u	������c)�32��_�8���`r�Y+����� $POO�Yd�y���7#�S��\��'U�n������e�T?�e��g�^2���ӡ�p�W�A�2��C�5H����n�	���H6��P����0���[�	��
�xڑ.=6�c�M����_vc|fAW��$�ϯζ{(�1o��z<�1�$S�ǃ��ƖG?3��+v-�dN�����=Z�W�J��(�||��p}�D��K5�nb�*&J�G֙ҽ	u��1H��<�Ć֕�Y
��T�Q���q����I�?	��3���rBh�z>�{�7�w�?DV'��� 2_Pa���狇��C�D񌰥���&���|�j�ߛ�Y�����E�^������t����w�^��k'���`�j9�_		�ݟj���vvkT���2F����AEH�g22p����ek�6K�ΐ�X!�ҼS�#La7�l;�����=0��횎���b��in'�OwQ��X�����v��]DA���P*�M�nWSN),(���~�����#w�SQ�S�0��yz.�w�~����^��k��?��,�r��CB�k'�� ��u���O�A�u�ǌ�IS`j�vbG��篘�����k2�Wӵ�1�:�2�k��א��̆84_ ��l��:�)#��;�J�ֈw�"�M댢#EΝb���O���l'�O&��T��P�"��@w-��W9+�
��F)��b���+���ϚF@���Bͷ����dk�~x��;�-K#t�$���!E��O�-��m��,��9<7��,��][�d>n��퓋��ծN��`���$%�_1�߂��re���1w	�}5��Ĝ��?(pI%��M��ZF���Hg� � �����),1bG��XW�y!��ˀ�����.�D
� :�o�;<6+�G�1f��z��&�{r��)Rh{����EYK)�q),�j
_V�9�^�����ɠ̼={!�[�F6�'_h�4:��tޑ�X����5�$9DySG�L�od��-�H#. v?>�)$���g�<>^+�������g��2�+����ҥ��N�� ��D�4U�*٠Rƅ��=��:� ����%���2�``��][?7��������yn�{�B�F��5�c'�=qFB�{�{�"M�3;�0��<R��0}�{�>o�=�,+
|�(+�"�����x$d���b��ĎyͦZPT����s�O>/U�eYO�g>��j��P��V��"��q��XA����|-�S���ٸg�;�!����vmh���ҡߺR6(�������U�
��PӓaD)�r ʖ<��Os�Ns�Y"��YX��ZXRi�.���laP��)GE����(�.�=ӯ\謀����9��q>��b˧tO�*G$5�
����5�J�ٌ� o3��|���lQ:�5>IvW�(-s�C����	��g�8�Й�Po�N�y�S�g3�k�'����#2���ġ
�[�h�\l��XSS ��Q������ڪ����y��D��ݡ@�fp�D����#ɡ`in��zc�cc;H�#�9.�� 
��#ړ���)�P���A�s�׋n$�b������%SS�;Y������V�z��)3:�~^gSu�en�:�ݯ��o�Z4�J��< �ǳ�[.���|F��H�{;����Ɠ�E��ncV����ϛ��K�{k�e���t_����Ւ�
��`��ľ�esJ�r�T$n�� 3���R��.^Ƈ��R#���_��]Ou�)�Ξ�!���gَ��_((�r���=eT� )؏J)�z������d�r@)%�r�B<V�vKlLU�怞 �Ob�����IjH�{���V��~�4��s�=6B��'"�W�Q`�j�!��r�Y�n�O�=�ب4��!=zt��q�� �`*���i'7��a��S����頊�������Nĺ�j�ݕ"w'8>/!A�O��vd���el�EW>~�������L������J9�ׅ㬈���+٩�oa0����BҸ(_;�}�+??B���^�ȩ�|Ş޿�x��G>��ȵT�ԫ��r�c���`?t��
{q&� ���艦���D�]ܐc
��O+�&ޮܐ�%qR$7!�{6�p�&&���Ⱦa�wTֶ�uک�<���H��XT2TNR:?�AW��R�o��̒��e�h����>��J�=J�%�W�2d!ϝ�˜f�ⲵ(���	w�Ĺ�o����� �<h�C�nL%e=��M]�@��Fm,uX?w�Q`]���i�����Kf��x\� ��,F�"��}�HJx�D����Ɓ�J��񎩆zh�b�;QuW<X���l+��qB�eަ�ÛmV؟��uT�3�K*)O�� �>��/��*A�F���&�.Q{[�u�E��K��~�/I|`2��� �i��W�*�F�|s����J~J�h�J�ߒX7�G"�m�)-�E�E�D6�+����t�;�)��Rt�r�7CG��Zݯ��@�+?��K"fr	�U�v�	��������+L���Lb�N�J�2����<�r�m6Ʈ���!3D�9s_�ZJ���"�k$�$�d�":� ����TǤP�z.gl�t��OS�ubR ku(f�;�j�E���\@��4 � ��ɗ b��� &��I����������k7�0#grܑ���	M����wSb�����a���8we��pS���<�8Ѝ�1���������WB �e��k,��"�̭(�rM��l��Lބk����6B`�O�ra���b'~�9Hp��<�b(s�k���Ɲ̌ڳ�`jm���1>��?mW"��0�:�9�޷M���BvP��b�+����
%�y�����!B�	���z�b�i?��V H��\�;�#l��0.g���o�`~|��Y�x�kB]q:='UoJ���髿��B��G����`��j���Mb�G^_�o��Ŏԩ�8`'F��k�����q�*�!u�5L�ث�o�D��d֤Y��;M����_gH�g�|c����}0$�<�A�t�eO��<X���/͸�g�i��� '�'��;�,
4f�z�������$��2�I��8dߤ�5�2�J�x��N]�s�E�H�ڿ��F0+^��\�,�<��z9��⺿����l�~l�X�A9	P��YƱ�G�KX��Ѕ���]~���NRS~c��n�N�.�zY�һi��a�U%#
~��u�H�����@բ���~}�N�QW�L��#||�p��3�T
ŀ1o���?�K]�h&���w�/�ݽ���a���TP��+D��������'�l��� o�(#jR�X�A����d�hf0����F�R�ck�U��=��,Jdg1��o�>������K<V������3�;?��EQ�?�u��F�
���A\A}3�$U�dDX���$PU��`�-&h�K��ӥy:Tc�c�Ƅ�:����̏�;�'�&����Ҽ9\b#��̽))!��5�_*C�N:����O�0�	x}��Eo[��w�j�Wm��v�n���
<��&���*���¦�!��K3^���-��	e�o��RN��+5��>F:��[����_az������Z�4.,���h�୦!��&M�����,0�r�na�Sg7\��6.����-��(�^i]��{�d���a��0���Q�p�"����9ZޙN@`Bq���T�=}�-�C^)�wo͖X�O���Áܳ;g�`�߃S�G���=F0�b���B5:*x��+�6��)����7x��F�r�!g O�m��a�AYƍsM(Q�T�\�D�D\hB��*��A��j�����I����z=�Ч��zFGڪ�H�ŴXf�u��@�S�e��P�U��(�S���|���b�nQj��Ԓ�U�����_��+�[5�7Կ�:�Ɩ�kT+�Y6
�s�]%#�k�߾B�:�^e�c׻5j�A�̥�*%"kQ;ݒ@d[��בՀ��R>�f�x��pZِ7�b�>a��©I1��ar�eR�'K8��lU���Ŝ�����e�2w����yB��nz4�v׾}��̄g�ebܑK��Jb��#M�@ЬI��<�0����*�c��"�(ʪ!��5{��+���8'|�����NPPH��w_�%�N��K�ز�?����X�(����ȍ$��o�(p/�bF2A=Bkd�ˑC$T���<P�}A�7��ʒ�6k`��ꖤ?�4+�s�h�a�zk_T��r�S��P �FE-�N�o��v䃕nFjS,�C:v��{��q���H��"F�4����v��蒽��2=��AYr�K�H���8�Q6�?�}���<�V4��ȡbT�S�)���s��#UlyJ�e�u�,R�Ȅ�*!�H6�1�����D�9����[����P�^���J� ��ǈ�ɱT�hB�zTA '�'J׷�;�s���h��/�e^����!0t�_D�e�pG��WA�0���� .�t�$e��oEWr��C�y�V>nZ����#XG�։�����e?�����8a�ޞ ]�7j�$Xbf��䒒9���].�FW��-�J>'d��{�����X�p�����AN��盍2����HV1��?w��z�%K��2�"�|
����R���G}��^(ZV�=��T8蒞�݀/�4�����}�F�Ă�d���j$+��N���i�Ĩ��
����ϊ����䓠��|l��z-���_���fJS���j�/��9�����&�c���f�6AP,>*��q#_�)Y���	��O��zMg�y�U���/J{'�D��^	�_it$�7Jn�>.�t�����k��d��Ф�,O"��v3�x�=`	�,W"�nNT��1��e�����Gez"qcS3)�%�O�3�dC<M��~���A��]&����>`B���q�Sͅ���H��jsH���VYQ����(��zJ���((���Dww����zh�������Ի?����;�C9�8t��<U��ǃ���4l��j���Q+�8����<�)ڃ�Gm ����ށOp:��m0�z�AZ��kl�n��<��dQ13SIȜ5C;~���V�h�Uyw���I���k��YLDsXs�A �b\��uu�H"��E��a��:�'��)����^���H\�e�xRe�x���eP�x����#&�y��	���$c'��@��
�^�L<���Z�W��9���SܓI���`��w�aԾBU[\�8{��XzW�O�o͔�4�I�+aԙ)W/�����c�+�D�7Y��s�h�K�i��f{.�n��Yy~3��7��+UB r$"�4 ��2蜁�rǆ���޺\u5����*��f.�1&�n�4�A�<(0V��$���L}�l����F�6�(�s`��mv3��#��!���?��{Hoi���[ԮE�LFg��rd8�W.l��4�$;0DNp��'�;�X'�J؍��y�ô$�%/���h�s��_ Ѷ@Z0�GX�O�b��+i�������Z�T��9�����!䆊��9���S�'�J$��5��e��?]l��p�KQ�U�ӆ���4�5JK�P�a:��Y��,'����O�>�p�5Eo�!�����cR:�x]sz�f��Ԅ ���߄�C|7����5�3��2�2���t��d������x��C=�ȴ��֣C%�0A}+�p��npj:z�:���K������WրO&؀��|������)�X���PȺ^͌V�t[6���'R������"5A��٣�W������_R�L��p�
�8��y�
��~��M��Fd�~�5�S��d3�6�EK<f���<V+��^��.da�ȩv4��Ԁުa���RQډ,c��-��~>����5.��iS������z����XdOSǖ�״���{�~���� 0[=c�\.�.��~i�S�ꁙ��>�{Z��^C�!�I�:��L<MX����Ys �A��dj,�j����kC fիq�Et������b�&Y$�R�ʪ��ۧ>sO�a!���CF��P8Q��ܿ$J�6�y}�[g��SG#@��^�ly�g�lz�4��ݡ܉�?�bt��d�=�*���8\�����
ϵ������¾h�J��7��j,�(D�q�1W����Wy�%���+�GJ�f�!�~E��
b�I7�!��D�y9J�'�2�ҧ������|rL6�tz3u�{-���o�}�g _M��V@w63K��vr.Q�vl�:����o��f��,�����Y�
���"#��N�F���D��w�OZS/,�3��-;��b�h�'e�3���#�C�D{oq;�c�PVf帞���[���m��,��yʩ;)A����0�^�|WE�1jm9ǵ�D�0:�\e;�c�����Ӹ1���$���7��Bx!K�.@(�3�B�'���KQ� �G���̤�;��暯�|cs� 3�NHl��!Į3����T`%�r[�cP� �X6�4�ڏH��"�%zm�r\nd�����M�ݔ\q��"�����ԍ�������(UVEgN�o��3���\�C��l5��qv���U�Y�#�N����l�n��ޏV)Zy%9�H���{!N"�^ .����ĵ�M�Z�焷��ma�+��hyϛ!J��̾ٽ�;����:{���馧���_��n�~G���!��"O�2��`��mV,�E�Π|H�#=g�%tIFz�rJ(�Gp��oG ��EՁ�R\R��n��ǟX�#Є��h�{��5Me9P}�ӂqA��-;�,+!ʱv[	����xv����.��Bs��*���	����Td6`t���	
�����]_&���6"or�����	�
�Y	�z?OL|�𦒪�e)�ډ�;�I��l�m7 #m  ��Kޗ�h��u%��&(�g2�S�ظ�138�L��;8��V$,@,%� nlz{�^ȍ�:�iUe�k���4�)�ئ�0 9����FJ&�S[BI�UAd���#�{Ć�;�d��X@�_�1�ct�q�>;��^ҫ3��L(߈L���zK�0���e���EH��M�Sr���,��e�n��X!�ꓽ�'N$o�o�a�!�{���˂gkL���P�L�
(�=�޳�f��ȳ�n����+@jQk�����C�#�c}I�9��M0E��ՇPb�H`���}�m\|k�Uc
5����\m�o~�v^YOWX�q2�ڛjNr������K-m���gk]�F�����b�j��@��EŲY�e��E��^j(��RR�b�f����R�c^P���c�6���%aĆH�9�,��`8#�Ⱦ\�MSҧ�H_�Wd��o���<�0�rmP�.�zW�1�x���D�:�V�ۙ�[K���s��?��OarR���B�ǝS��b'���	lK�ÅP">0�]��ˈ�Q�������H��ݕ�`3j�7r4#w��Ȁ+�J���O4�T��W�Ub��bc�*��?�u�\mΎ�2�@��ǯa_(ŵy����7�m�C/��i���~>�u7��<�}㭽����:P�N���O} 9̞�9yPq1�+>�1V
��[Gw��:/���)���n�4owl!�ұٳ>��#��?7Iޚ=�U���;�ء��͇��7d��w1;>aZ�b%�H�F�?#�n��B���:Ŕa�~��WP_�a���ഗ7����-٣A�|?-.:~Vb��/v��������))�g/����*�C����o�XY��|_�\�_c��M����Z��
0�=���Xk�9��|,'���u{�6�C��>�w��� c���=�}������4���������N�t��
��2�@��Q!O��e%�XӖ���J-Z����T�͇޿��I�#�wi��@<��Z���<M�,5�>9�,ݦ��y,����Di��Mg��a�C�kM�y�	����۩3����jziϳ-���ۂ����@��A�qÖ/��B�c�- [��;y��������"ֻ,_%$M�390�ހ���Q_�e��T��)�t�*ɀ��"�I��0�x�t�֪T�r�G e�d�!�u3��t�
�y���}�3k�5����$ �P]�����x��`S |����tK�U���4�a��Dه�OeE!�e*���f�JlȤt]�AS�lAY����ᐥ0�K��'o]��ɭ$D�zG���<I��U�������*b&~��vv��h(߷#ak����n��XTz�w F`<�er���ʍ�.?��3F��A���c�{y��W�H~�d���!���A���w����,���-�UxOY�-AT[���э؄ _�k��ܥ���z,���l�5
�Ci���PK;D��z~�=C�7=�y+<O��rv|�#4��PI�8vd��i+b����~��q�ϭ��޸�PH}�C0���	D��{(�r:�u����$�-:���(�*��m�YکP��C�j!r�!�[��У`�(�]�#�ŷ�c����'�!�B.�t�j(�B{�[~����٫n�B��Sʁ�U�����	�X�����%�)� �"���OF��Ba�7���~��&�*ؓ	o&vmW���IRE�z��њ4l�<������
7%Z'n.E��{���JE�FFk:V=�#(����H���5�� ��0_ٷR�l����=����Uq�vo�*5��Dw^�F|���&#@���=A����V`�ˉ?���<@����:�/M�Tkg�:�0��2y�̶�62�u�AeDM�֋���'v)�`l��{�o����Z}$�P�`��WbA(�: ��-�l����վ�X�r������i�Y���A�U%�40�wf+��T� g� J���B\򖋹��@v�#} _�̊����5T�[d��ַ�x/���������N��ף�Gf�~�L�с�6no�)�D�x]"@�1K���Ʒ�����G�J�i����~� � �)y�����wt��j��6,(~��6����q]��D�Uv!�M&�	SԄ��>������ϐ��/֊9�7dPNB��x�yX{�K)�`�(C&�����"��ұ�ԗx4h���{K�`�;������ S��)��\(а]`�h��kc55m�47��,B�C�3�e���s�b���O��&��ތ� ��W�� ]G�豒�/V'�,��,
���ᙼmE��T�jN7,B�4@ި��d�I�#9��g���e�C��f~- &�.��h��3Ѡ��s$�
����l�0�Q�ƙ�4��q"<G1w�=#J$����w�����3 x� K5�]wZI;[��_@"��=,CI�w2�Φ����35��݆V��6�jc����)YP)	C��B���C1���w��@�����v�(��h�}T�Y@.?
/߾E��(�:���Z5����x��Ԑ�	sVr��^���̸ӻ"�_�E/�����v�P��EN�q%��I�\�$���H��Jtj�6�$�Bv�F���)��V]c��;�|�v4��C�Юr�q�mJ�!biZ�{�-��CDϜ�P�
�������9r�Ml��y��M�W�����^�K���� ��˾�������?���h^���L��b~���!�bH9�\Bn#p��~���_�F�%�����Qf���z�n��ZT�v�����z�����T����]�%�:���U�W����VbН2���g�����t>V'��̄������@2B�t����ˆ�1�k{�ȘLn��
@f(u�U7���N���J`�R�D�/Q�Y�������f�v�`H�H<�k�JY��z�z+�}�3IB�z�c���tE�ܚ_q޺��G�@��gE`�ho�,+ۗ��y���>X>�٠�����%�ѣ��gD�e����q`rG0ذ�'1��V^�MJ��X�Ӯ���<� ����+4�)1E��A:�7��]�6���)�R�j��!�]�L�?��>;��[��(B�y���?bVA�5\I�8�&<l;"���R8ôuo��^*^ds(��T�������`Hr	bu�ԑ�@�Y��
y�F&5	5ܷ�ϜL���(�Ѡ� ~z�����͔��2j�<��o8����5 ;�����~n�/����G��f�֦�f���ӉS�s�w\a����k�lOI1���;dy%$����m���� :�oV�䇩0��R��T��?��B�ԣ��-��(%-{Z�q�o> �K�+n�oql��V�t����I�� >o��E\�Wp�.���3�=�悝���/���C�cV�
�)!)US��=�a�x�o%�F9/0�x�I)�)�&�y�uH6�QZd�1{b�N0_����7�C��N��ɧ��N����6U�0�ay�40*�]G���ۣHD�mR���Ё�
�ֱ�����2���h���l�H��K�E�R
J'!��+���@�j�o=�Q�C	�V��y�Y�*O�������c]��%L�քM�����3��w݉��T�f >�W��~�p�\�Nc�=��q(��z��]�*Q����b�di�{�0�ı�FZ�f#�����Ml-�æܰ$kFK���2LE��.��Y���5�xH�ì�&
�N7��+��}nSf.��kK3��/���IsTk��6�(|!��j�%��"��x���;�r�ѕ���P����M��y5Tz4;�aE�$���g@���1JnvIpi��"��-�n�Ѧ|�-����3�H��r�aƙ���f��O������5�hL&�FCo+T  ��A[l���)ƪ����UK�~�u�����}K� �_�M�p="һH6��/���_��V9����G�}��T�)B���!8y� J���Ϙ�6���&���.P$�dM��.�UY��G���:��(�C���?������T.ߊ���V��yu�N�:��m���OW�)hm��pGOv���C�µ�pM�-�ϙ(�r�W+J�M{%TWEC�O��@F-Ī��ò1M�1i�r �*�~ �'�� Y���U����Z$m(�k��)H�oM�w����Dl����Vo���� /��`�Ӭ�!�M]�s{'�蕸x�U���	��x�n>B�q���[#���i��:���/��J���s0����
~�OК�>��e��_�TJ�S]�e��oJ5;����ac%�XE�]Yx��?]YڿŊ�.�;.I���>W�AlZy�l�����}�B;3�B������ȩ�>̀�z[+��������ɡ����3���j�t@E�O4���hd��Xy����"�啢`"*�$Q�:��S��i!y3�i�s�xMLs�+)�۷�ζ7�;�K���
�)�����!h���
�*s$U����E��~�[�ݬo��}����=>>/�:��S�0&�����o� ��^a8�$�x��nӫ����]�U����;�鞛�Z?����e�wR�_�ob��5�ߔ�e�\�4�Դ!Q/�B���0W�V��5�۵��E�тO0�	E��=;�n8��%���w�7x1��0�;{�o��]���% �.��+��Qn7���u쮛��/iJ.q��s,�~�8X��F���(��רU0�<��y���P�vuOtUr��~�ǩ{��f/4� ����!��0�+{���o�`qǶ�v��- %dx��_�_��*c�u������7$hK�M��a;��
U/��@0cV�ȰZ4@����bk���C"����L�?��I������r�2u��uр��D�(���x�m"����'��_�f3�؏0��D.Ҭ��=J��8�m�x���c~�խKU�=�~��u�#e�FURg݉��|jÿ	x22j�<������'�P�e'c�(���c!��	���iL��C��ʈ�hbN���?��v�H� �\zZ!�-s�!�p�!j���>zIct�7G4���	�����p�B�:���1J��S����Hx�i���qD`�;�!�;)�g�wQ�
g��+�O����ojS���L�|���~��'@�\.��
)u�E��q���'�rW��3#0	eW��h�o��͉�x�٘!_`#ԗn�rJП�N+�c^RsD��ۓ*K<���}POk�P�W��)-�+L��Ng.��FU�4����O>��s��]�G����u�ؚu����#��c ���U����+����,^u��u��Bni��P�7�1#���9�7�OPET�@�
#��7,F.��]��'��E�~r��^w\�WV�a4|�)�����t�?*4�i�wHl��-Hv)]�qH���3�d%W� �&���ry�����W��5�y�p�mw}�O�;�@k���X`�|a�oA&���)��KY�#��y�y��<$�����P�vܔ�T6j�_�e��sq��u���o��#j����(�i�?��+p�>�8�1��7.�ɭ�%U<�h)(�T�y���Ûʲ�h��&�l�#�݆���G3OƤ;�b�g��Q���.1��3�C������b�}glQ��C��v�����3�����r�pTM���	�݆L�]逜�x6��u�En���PY�.���z�,S�N(A�I7���M�ͫi�6�ۙ��ļe��̸�Ab	�Ӧf7�W�7�H��T,!����w��;��d%o���b�E�?���-L+\0�O`���0`B
��ˢ�23������}}~K���ⰻ���}�K��현N���ƨ�D��nR�fó)=^��~*��BP��A�5$
F�;��s�fnVZ�ꠕȪQˋ{�O�EB:n���O^�_5�N��p�C�`#Lx ���X��w��E9b�ޮW��L�����i\ǩ9��3����$Q�
���OA���]��'\�E9L '=jN�� Ʒd" �>/��B��z�T�Z��"NЧ�zAJ޲�6�/
����οcg���t.� �]ㄅ�7�3����Ő
[�H�/Me��*^-N�,�֊��ИP�2�x�͈��1bTr��.��8i�@�K�m�B!���Sv¼A�O�w1�Q�$�]b��&w���)�B&�H,�p�	"t�iC!N0a�Xݨ����-)���[u�s����5�o'��VK��<#�t����&�,D+�<��HNg�g��(��-ar���i�竜w�/m�z��6ӌ��a}Aa��*�9H!y�]��40�lw� Q�B��**�mh�� ��ΐ�f-K�Aњ�x�N�p~�8���duK8Pf�]��.�F[�$��u��Ь�\��Z��Q�A���.�3�\o�X���̤�d{����,T��J��G�_4�J{,�H �2i�1q�=Ds�=�u�̦2�p�:蕶XǋB��7��Mg!"�;D!z���6�����7�|��c�J�H�2Kih�@���+:�G��A1P���$�A��<&-����i��,��d�D����&�R�J�2�8���?��#�=���!�-%����v��P�-���y�m8#6���Ns8y����M�27j���2�a33���;���� �&p{��4����gLU''k�G2�[��q��2��8A�q'������-mH'i�K�gs��=��{�wZtF^���[��gV��?����F��ˈs��������`�ȂKDt�:�����AЉ�Iɹ��^��$t�Tmjm�i��{�}ك�?Rq��7!?ۧ��^|��Қ�̚<��rw���ΜH=���1a·Ѥ��ǣ^hZ�RN��X�O���yt�w�L.��y�˨�BX׮�R�~ί�ނٿ�V޲ �0��.��(U+�X7Y�Sv7*��q�ɗ�ڱ��'��x�7-㷱��7Lx4)�����ݯz<+�g��s�C�;��Ȟ7>���`b�Z:��w�T�}�Ú�O1/��
��4��*�X�Ϧ����A�?0"��K�����[���(����51{�k^ק����1���̪	�㟥�������.Ӆ;Y��z�/���˚)�>�s?#�M��z�=^RMq��v����ZT��-cҁ�*D��{H�LH�xZ*��ZV�R��.F�͐'�f�Is-^�~ސ0y�zJ���ֳ�^A��I�Z�{�y?o%�(��B#.�.:^�m�#�pߡٞ�[�y��۲W���U��~��r����<��Cl�q�����C�X�o��/�|I �?=(���B��78e� ��]�;�*ɓG�(��Zt�sw5^��^�_Kxs�`�]�3���_�M�/L)e0��H�}��g%���� �������ENS�%;ױ#��I�`܊f��Y�E狠�qF��e��1�ʏ��?�r���\B��p�ɷQ��B��i���x���"���=	ВzV�5�&�N#��X���+_��	�����u��?�~;ϒ�Ǳwk�~7u�ݦ�<���I԰PHZe�4��7]�+6TB6�*���j ��R�I��΍�S�M���6aAv�X�0��s�'t	9�A�/6��� �r^��q�z�b?
{=J��M�ܸ��1+]_��"�f�|#z��C\�(A�eE�tDܞ�����"�j"*��x9n쫴����hI�YM��y�8)�;KK�|���"�N��R�Kd��A�u�&#��+<!<�bO}%�*��q�1�&bz��!,a��������Q	�&�,��X�Į�B;8g�P��Y�և�
��֊p5��̘s�خ��R����B&��
I達$�y;?l��׊�Ǚ�5�+��Z�K�����ch#.�r
�ڄ��Z�MW,@$�-��)�}"}H��:�#]i��ٌ���d99̴�Y����n��{��R �Y�o�ϒ�6�Fdo#2�s��ٽe#[��\
������!�Z�=��e:�"ʟujX�礒��N�w���n�x��DE�a�Z��<rZC��-f<0��v�4}/6���;���?��V�z#a#NAk@L��Gn/�?]Ϟ���@�'�4'�AIY����͚VB�B��i��B,F���a���Fu
���_;�~�K��٪T�p�g�t�<7���A����WN�ʷ�g�]���̲�9oZ�N�X�nn������3�?+ٶ���o�~�Б���<j뾠]!%�6R�y��´�w?�h�x��gM۝�ݦUF���`�T�MN�����f��;S�	%f&���b�z=7�+�x�=b�ӟF諐�O!���w)Q�*��}[�o�� �W���Sp��S/��3��1�M_�1����B�U�#�5Kk�l�Cς&s�{c���L����aO[��*�"z�j0�S���ff!v��	���5���[�v�W..//kKY�]>��Tђ	�gB�//�������-ǣ���cu> �k�[�O��4�+$��*׺�I!ZYdXw£uf�8�e�|�kk�z~3�B�hI�o�r��w�[䷼�����t��X��������w)`$�T�ŏϤ2T���O�u@�z�]�	<���e��d*��ȡ5,k��Rl9H��V����S��%-�+^�4፧�aO;Fa#,��o>�_���˻cxi�o (�Ӹylw�B�	��h"ʀ��+�����An�M/�Mu��^���RX�T��s��Ϸ��|��Ua�v~���Qר���~2N[�g��R4^��q$Xy���2��m�
WGKv}#�����-�������y��gb7 �:�.|q���1�&+�W�f�>oP��(vu�O�÷���"!}��;]��"Q����#�S��s�p�����ʷ����C�߇��?��?>��*��'���\ �ƃC����N���I4��)�lk`*o"��a����v��1�+���иR��kkd�:vo�����6
�o�����UMc��'�뱦<�ʿ�^��/�Z4��^F������R�s�k*�ŎYx�~��LX9���;�����e6#���@eˠӪ\�h$�����
Wk��*�sj`�,�ޠ���jFP6��zB��#[/jn]h�G�&�57��ԭ��ؒ���X���e�PTB��6�x���-JH��Pw���H��{0��j��󼈡���w��Ab4G���ɢZu�����,uJ:��� �T��3���sA�<	���w�1���HM��'���Ѓ�[�8H')���Q,.E1z����6}g8��rH�}�i��_0D��T�+�h���z�X�7G��Cm&�O��ӹKgT���-#w�8Ya3lQ��v=���T����ߍu��xv��q��	�UX�[���KO�u�y:�g�l� �+����]��:����+������p��)<����Ph���Яł�5$����@m!���p��7��B�˦ű�b�X*�OW�_f�<.���8d:�
(K���έJG�XK|�u���^"�[~7:�N�PȀAu�.���Q�+[L�ây��	C�����`;I���((^����(X��	K��0P�_)1@��v���P�<4�m~�f�+Rs�9�� �.�uY��or	����R��n�{^Ҁ˫ҧ��T$�H+ݥM���y�qD�E������5X��*ּO�Fl��,�/ͷq��Hm�}M�ނ�w��OC����t����8b����3͒�OQ���~���bļ�xj���umN*Y�����<z��s0qq ��v�Mپ���|ץOV���h��A�lO�����+�*Z��^D:��&aG����D���[1�]������VHbP>�9�E64�����
��z��?��p�<2�Sc�P�[խE��d�M����)r(�#� ������s߿��m2#:��a����U8�@Y�&���VX2+
䬻q��z^��r�L}��!ج}'�d�q�^l$4�1bڏv���kB��*�+���������g�T_Q��f�듮�S�[xJ%���<N�z�]#_ hn��a��JH�)/i�)�*�����}	��^5���{��6�"��IC�;ٹn���8fI�OȈ���4X�*A�����;	Wmy���6��^���x��6��W�1���iI�_�Xcz�6��ZBL4�F����!������"F�n�?�#����_��i��/�D;��g0%"{��W��4x�PZa���I�̯��s�s��h�4
̗\�AF�i`)�-q8�����1�;oZRKs�~PW���1rM�B�*6����'����^{�zY��h��Z&Q�
!sFWgޤg��^��)��1=
�kd��V'K�QM~���j�\�9����^w�&����s�[��f��2(|x�m��_��y�{�˽-��R|�~�Ӟ1%g�(�������N=q	8m7>���5��Xy�Ў����S`�B������K߲���������1kJ'C��e����^�"νd��D����[`��x�BGv�rCBӝR�;r;��M�
�&�p�499!&�`�EG���[D�ڿ86�(��Gz̩�A������!aO��T�ʅ溞���i����t�٨b�d��(�yy�}K)�g��+���Q�p��5�{�^+�J���>:t2��`�m@$= �����Wkt@�n�2���(^��J#�q9����VV%���CB�Z}B*�\"���3�I�&� ڳV�R��ל�܅ v[�66�I�h�N.�6nɢ���������~�$�o�T��#��h�֤NPjwo��Ś!����U�B�|�:��n�+�GI�)�b!c�M#4�?����);6Wl��\Zo��
'��Y�K�VaI�^�es=�����Jϭ�������d����`-L������캝����X}���.-��I5�
n�7� c�s��u�@Ӊ��p�7ͫ��FM�T����Hн�){���il���t���90e�Y<��^^N��v�P[��PE�߹Z�1檅��$�qܙ$/N��O�d����6!�O�=�>&ג��1E�+T1�iO��n�aEΖ��m��Ie�kF���T�{G2r�uy�����.���GcJ���ݖ�-�!�<�����D���.0>j&����m�H�$�8l�<N ���Հ� ���U��6��Jڒ1E"&����߲�~+D�!���g�q����56�Z�utՌ�� 3w��r��4��mPc�si�%J���;�!��p���C��P�r����������ޗ���g�U�q0�+0>V�|���"B8/����!��.�q�p�^+�e�w���N[�E�i	V�iC#]�h��'uh{�K��L	�ZN��O�T� �]�	�W���i�mw�o���~�3ݍ�	��v�$���V�������+�No�(���&b�%���G>!)l�'.,Ȼ_�nx���z�1���|�'��@(��2M�z-L�4^�ޟ�%�]��r�Q�*nr?�a�+�����1"��]$��_�=�=_��:(�pD�&� ��L��E�z�4�
a[>Y�FͶ��sM�`��aXw�s�� Z��ԅ����M(6��X?��@�Zk�<!~ٙ׍F��@2�;s%�YҐE�"�&��"�F��lR��(Lk�L�O�M�j�$	�o������Zi�S��+��`��<��`�oR]W~�������
�[3Y_`��|�o!��&|i�y�O�*����>�eV�
�����f�*���ŊQN�wkHu5�=�qF<�2��EPހ�}|A�oI4���C9
D1���J�S�/�E��h�fW�~����Lc���@֙��ũtL'\�?��g���e|x�@GPR<9qd��Z��ZW�	��=�*�a��8mK�n\ YJ����f�(�P��o��LjJ�m?���9�7`�q��ф��i�׆���W;����R��o_^�������h�*�]�&$cF���FU��n.�|
͜��/�����I�����Q@�������8�S��>�{���&�z�CS`b��^P��n�W�J�Ϩ�6d6%@[�$�|r_��ѐ���i�N�*�#i�h�\	���
�՞J3�ޥ�k5S� ��9j>aZ&��D��Z���G��'D�Y�rǵU���`B3�j�5HW��nI����u�G�A���:�}�����9U$Z ��dДnb���<�1���##QH���Q}�/�Lm�=�а�A X��P�!���&�����]�ۋ���lRz�$���IH�fh�d�c�$�&�\��~zN�'���9-�K���n
"
 �h4y�B���͆4�Դ�T���VlZ��0R�	H�Uz�͵����zq6Nmݛ�#P����2�(��M��dz��ɽ��z�������#�Y5���4����q�7����P@�pQ,��%�	y'1���a�wu]l_ a ,7��$���#�[̇ V'~H�`�ٸ���.=�zp�«���0y�/�1�<X*�B���#
�;^��}���B���I��Һ�0e�6!_^i�&l�53��]�+k�s?E[�O���9-oC���j��Dw�,�[�#N�L��8p	r����DS���M���.�4x򣔩Pm�;�D�<�
���@W��d&����"-������$0+(7Va-lO�/.�@]�d�����ЗJ�h���7�\��!�5oV�I�����{����ѓ���s>\9�w���S����PvST��o�T̼P��}�$I�1��@��(�#�G������;sk�;����6Q=����:g��/IK�!�r����g�5n���.B+�/���,��u���X����?cKX:o�48X2�	&�U��I��C6��1b�g�~*��@ �^��)��
���϶@K��F�F�x�X�c����&�����8�b��#�H����{h��FQ^��W��#�c�p���̡�M�Z��>upw���$۶���y�uL�KC��aa�Q���3\&Ӗ��� �8��ɠ��L �D�L�kWY)2�`�'9�}�^����MY� *�o�j��Uo�%"��w��ϓ�V�Å:���E����e\���_�������k��OƜ��:`kN��/�u�mJ�X�V�p�6{� ܋�^R���9�'�G�A	 ��3�#����o��xe���<C=/ڰn�)C� �b���|z&���q��	�t	Y��/�s7>3�0#0����A��H�
��ڪ��u+2zC~58����.쑚ݜ
+�\	���'����3�>��IL��D�����: �2ՙ 3�j�`+jϲ��?�ɮ�a����![c�v��?�< ���ZI&��g���킏3��I U]�,p��/8ۥ�vV�=��)��0Ì�A�O�=u�wa���\+�*�G�t`���GA��I�Q܁��-̶ xp�6긌�L��Q�������]���H$���Rrg��zW����n�%m��?���6D�i���c�lǦF ��,Of���%a��2�	R"�s.�����6"���t8H�,KO��ۿIB�Κխ�t��ӊa<�� ��E��5g#".l-rQ0��m���ܰO�;��n�`�\	#�D�F�O��x;�q��VG������tY�z��3�MA�P3-��w���ܥ@�����Sm�tOMy<xY��[�fT�M�e?�̠&:�P�'7�]
�/!6�S��d�һu.W\%�m�*����,�2�(�>+-�P��y���i8]�5<U�^�]�/b���\�Ɗ��U^��_&�>8!J�I$3��sRD���S %[y;e�_&�����%��9��|��&g�9L'\�!�����[�8����ua��Q��Sd��9:D��xp�6�
�0�E�Z0���-��k�o��W��5h.�'0��R��V�f�
�s��u z�Bpl/�4���jf���k�e�'�%7!�u̽n!Iҥ�^�zf*H.�vVo\F�Or�i4�����m���^�#�߅�Σ�d��PL/�L|-r�9�f�5�7��B2���k4� ���il�|���.�U(7�3���0M��&;���G}Q%@2���6�.�AjJ�ݚw6�`v1(��[ya6�l�����z�W'��j�D<���`�)~��Vm�#�f����U�N����Ch��a�ἠ��/�݁�E�rH��̑Y��4�� ���
ʒ�����@��t4&%ce9#�7l�"�7����h�|�*w�j�d�'C2�#�m(��k��]�.�0Wf�$2;\ jG��j�u�Bh�R_�!`�ԟD��R�������̂6T"��}Y�9��� �<!���͓ !���jȵ�_�H˙�d+��A��F��U�XCP�+�K���ۙ����X�Q5��|�y�}l)3�k��_,��ǆW�;��,������ {d��7�� �d�V�>��b��*Y�����0C',�4gH�ϳ��Ak�pBK��	R��D�f�h��%Z�w��i4E\��q"D����#�����S�๋�zi+��EI@rN��:��X��g�,�/܌��Ʋ�� ̻*/������N#�( �ۖ@��6�#j�Wm�̃q��x�;��+P/X[u�g��2�,!�6�|,� و�%T�q�OAf�r�$�ds8��C,���J�<t6c�>:
�][=��'n%��%���#&{P=������`�c8�E�˾�2�� ��{pXU!֢,���
�Z��:�w�\8~	�V���W�lh��({E;��LccC�=�����碲�$U��UX��qK�+�D���"���� ��8�P�"i�7xP|������R}�8��F�U� �����G���9��זt���7����
��B����s���~o���'�7�,k\��es��bP�Ώ̿1����o�Pc����7�0[\���~u�0��"x �TW-��ٴ��g\��J��K,+���S�Rl��j5�m�!sl葙�@e�,��T��D�p�5`�Mkcڂ�ˊ����E|#��� 	͞y���=)�nM+~� �}��:hp���%�"H�ڹ*RZ3����|v"��U�����Z6�-����$�Ė�[�PyvOy�{��.��nK��"�Eo����汲���m/��p��ec&�ofZ~���ݣ����������0f�:������M��/m~�@���(�u�ƫ��"St-e�h�Tz�-��̓>Q^�W�k�eS�������T���\���uY��P;�i'S���C�W�C�du>�{t���\+۴H�t�Ř��͌.�~Z��ަ��S�+��� �t'�{0�O��w���@<�O���5$A��8�bJb���q'~�,(� ��4A��-�T��~���'z]\©�����֟�+�L�5C��l�糭%�H���A�m�0�����̛����&jP�`��O�ˋ0�lf΋��)�mt���"*f�|?g�H��k���YfSN���$v�M8�E� �%�����g�.
��!�	��. �w��\����2�4N���t{�κeD.�a��݊1��c4�*«�Z/�}n8a�<w�f���*�cT���*�"�/O��f�E>[����	w˷R�����]�`� �h���
c�MRF�!��v4+h�8YT3fs��t������4d�(�y��ֺ֎� ]�'�LVc�B97��{��5���\���9�b5$�)���Î��$��u�l_K��Ede匇�Su"��}��<y���&��c�#��<��R�j��[�/!x��F�1iaxD<]Ž��WY����y�:1 (��\�x��
����V���oR��>F*���/���Q2���� c�2I=?A��6
�:��U��ɰ~�=�m��`�����+�����0� �sa�����4�f��I6�\�U��3C8$�YWk�����^�A�������X��/�z0�zK��$�@�|�1}W~�����$Yqdco���]�Ma�!���Ra�������;9����5�����U��j�2^=3�@�k��՗qH�s5f�P-R���ߨ\:�b�^������`�15e���*���Fbv��/�9�4_6`�B���[��a��q@����XG��Z��(�1�C���y�%��\~/E���Zگ��?;��(�[�_��p����h����t]ͨ�d@�BA=L`"�A7�0�i����~��L��8PoɧI������S����lw��l�۸���>����>W�M��M爑�N~h�J�lXЭ�K�c���ƚ4�W:�m=a1}-�vP��T��&���y��6axysG��V��tXѫ�e"4F�)�ن$��A���8}8+�S���R�D�����ȫ;n/���(�G�dޏMYٜ�.u���Mt�\�z��W��jV�o+!	�ܥ��z���+e��Y���s��nդ3 ��Ugp �|�K��!�y���p��a�J� �^��b*8���L�PϯsM��Y��8o뇠L�`Je,����:G�E���]<_�Բt�R�٥5#�DR���S��*��:&?
��,?��������+��|]Kpqz�2ZT�Ҙ0�3�☀o©�>*�a���*�� �%���e�hԪ�	��-cʥ��x����T�C˜�j�d�ע��b�I� �l�M�r����}�z�|�{�wO�����2���-�����׾�7�e�&�����:?����`)��U����c8/�zǗ�M7�S~b3�z.��Wұ�Vdi3�Te�|tW�Ӎ* `��E���L��wF�V��B)��0=!��Srvv:6V|�>Hb ���ѿ`��3'ql���(�鋠�}X6���8�3uy/<�>1��ލ���pF�q�b<W�eK�����KB�j�=��|;hL�f/��q�����nV����ro�bɌ��3L�>홞�C*ϱ�9�g�x���ܠ���ջ���Jq��Q+�siy��7��Ι��[V�_�EGw��{̋��m���?{?47d�G�\ET�(�d���?��__���^h���H��1�B+hU; �5V�"��ńJڨ��By�~Rl �fw�H�X8I��Ej(�{��m�_�8u)yl>2�G��	���5��rh�;�(~�G�q�<mb������� 5c=��oC\���F�̨�Nkk�=��VY!��Y�UC�8����+���;ޭ�a�l.�8̀��ͬ0+Vő�@V�"��Z��Hō�i�J{�����7�2�VV��%�����@�i�ܢ���6
�e½2�����$a+��_���ЕGG���c�����^K�O�ɰ1<N�Aw�NA�7u+�8NcR��,r@l��b���߽�G1$�ĳ��i�H��<��e�(���ADu�����i�9G>7�[����V�)L���q�=�t�}� 4ĝ��E����f>�UZE�L���:;��#\��#B
��Z$����L�-����Q���pN�z�;s���M�IP�ؿ���o�N�Ζn�Η1@}J���*�v��ŗ-pB�=J�֜KB�E�XT�7z��3ɢs��J�ધa�V�0������y���/��?L9�6|����"�de�_�"ڌ�ח0tܶ.$rhc�B��l
I~���"(�?eh��1�p����^�l�Ƹo�藺�l�o�tyh��X�مĩL��aɟ��ԛ}��AۅO��6��:&�E�6l=ޘ�w�
��Om�F C=˸N��q#S'��o�-	j'�?����z�3�k�8��~�L�CF�%����	c:�!=��\���J�TH��q��mK��r��Do�͊]��籑M\3�1��&�!�����,@���#�dEh��R
wRA_���7lq�ʈa��.ӫ!Jb�hAh[O�$���Bg:��1-�s����U$`bs1:�䡽���7۞����^쯊�����W$��&�w>�|��:�%#>R��`۪�֚�]�!9��������������. y�@����4vۧ<sI��A��l՜B+�Ϛ�ѝ-ٗ�����h��L��9�H�v̍��?֯�,j*��K��rbҧ�`r�t��N�b"��s+W�����O�+��@2�/M{Ov�x�� 3+X�"3CҀ7�d�<+h��m�����߉[��+�;�����=Q�e% ��Z�����i[�W"1��ͥZ�8sy�P�}C4�>֨_�a���#�ĬG�x�5 J�%��0�1۾�ўG��^�^_�^��P�t�ga����J����]|���x]7�h8�り{6�!�c\�6��6�:�rW�k��_����J$��Oo�e3!��7;^�$���0�I�2�KGX>w6h�Y���#j��B] s�1���
��m����$��)�����Jwԩr+�- �߈�;� �ѼK��Iƌ����Mb���C�����B���܆���	��a*.[	U�@���yf�q2�9��-1g��=}}	��	y�s�Qy4�@_�Q�
ŉx�l����	�K���7ك�7o��r�5ʓ��x��
�
ȯ�xlG�h��(����y�����G��E��X�s�����LU�<�]s���K��^�L+����;�zԽ�<�k���|��2[��i���QV�#�����_�k�|�j��#�lQq�F�D_����*�j쓡��a�8TڭpA)-��z��%�:k���LQu�C#'�I�j��$���X���g�����g���%Hyÿo�B����q�6���9w�Z�3�m?�?Yy|`SѡA�T� ��Fk���# �-���� h�@���9��8���!o�������Me?9"P��'��5�E�g�ߊ�ۤxS����Yk!P��8�&r%J�/$�	���s!N��1(�����Q�|���uD�(bj0��d!�"^@!.�X���uf}�dxme�#�K�~����P�H�j�;�`Y�3#kQ����9�s'C� A����4z�V�xg�hX�1���gc��4"���ңV�,�������moxm�����,�Οo�ޔ��=9�9�( %�ـ^�D�����L�ݘ[чSyabz ;^��h��n���P��H� Л0VT�_�{��=.�FA�=��S5fY�hr������'z�~�W���^�w-"m2l+=�K6�s�fͯV�� �Oo��ʇ��',_���}�o��R�q��*���d��+~�/�,�Q�����C��[=/��I��u��Q��� V��v��-c�kɬ�x2&��9X��h�����H<�Œ^5n]�A�D�M
�9�i���Knk�77����F ��`TVIC��8�:�)q�8���!���b!�l����Y_\N�T�E�|�.�q���+�V�K�_�Z��Z�*���
1�g~�_�0��)M�����%������!���$�G^ʏ΄�yb��v�À�p�t1���B��~T�bQ(Zݸ9� ]��ރ�b����!r�O+M8���������P�X�&����.�%=9!�Td���jÚ� V��5��ie��6��8d�~ ��xJ.���u�D�-1�F�"`�����cp�GCo)�ݲP��>��~$v���;��ef�=��M���qOfu�N��V�.���y�=R�7k�qؓ�z䫊8�j��jbb8I�n5�_�/G�Ⱥ��<5�7[�:;����\It�4K���)iv��-��P�u�{��[o��oY�WE�� ��E@KN�*�@9���c&�������מŮ��D��J�O��/`7P6B;Dr�JԶ�+�,]�7�,�S���W��V�I7�P���0�U�I�|X8F<��P�[9b}~�B[�G!'vB���c ���dܙ;e6N'���Q���=�/��Y�F=���p�!$Gu �in
X���m�s�M��oe�w��b�"���C��mmG�g0�|x��N ;���z�ʌ�����Xm�^/�v�el�u��
`�ק^���˓�]���6�I���}i- �1"��m ��6at��]���V�zR��p$Y�<WX�~&���Qo�HX=�U�k<�O�ivw�
̘�ĭ�{�;��Ń&10o�j>��+vU�zE�n��yc�0Q����_���ڔo>mM�z��}�+�䂖��'].�!��	��P��EE���������]�@K��`l��UM��=�����n��nJ���>7���3�e�&�Y5c�sߜ�N��	r���f�F�"m��#����	��=p��b={�Y��FٲM��4K��ˀ���?�@������4�{�څ-� ��{pi��=�a�����3�)��(e8+�ᣌ�;�ւ�'V��g�[J��Ml�u�7�#D��P{UW 4/3�^ʻ����ݤk����K{����luʘwY�)�P�I+�hɓ !iԎY/���������W=p8φ�N�y3}�����n�&Z�^�L*�j3��*�M�^U-�~)م�k�6@��de��3��QbO��k��v=���:;�%�s�|������!9
���Y�]6/
{��q�(>�D��V�ҧW:���U�pXNc)�Xn������h�$xy�F�k"��"��(+ʗ B]9�q��>�J)0tm�.��L��P�bѶ�^vPゖ�:Q�����ñb����S-��+��_@�R�P�$��Z�g�B�JWͳddd�������v���-�z}���8��D�vZ��E6m�~x3W���(�*\Sb����A�EI���\=�\=U��o��i/}����8�D�p=~$��	lX�1Q-�z���Q6E_��'Yk�1��M�ǻ�i-�j,�c�	�<�g¬M-�(Q�������w�0u饕���\eA��@(R��8����A��z��U���x�)91�r�`?����3�2��� ��.�����ђ(Wu;A�4#+���}���\���� a<��p�{z��v?a������LOr�uΊ )�[��*Nl���R�3јe�գTL&�G?Z�ьM����FT���ku>�|��f��8A��]������o�+3
Yy̥=�.��h��g2�mj=�t&i4cz�4�-�/���R�A���Q��ܝ;��L+h�ü���?�b�gt�E�T ��{u�4�:����Q��	Rͅ���YB�D�67���Q�F�C�i��<?Kj|�d�uȍ�==2RP�����ۻVI�QIQ��bdX��.�5�
ݸ�m�l C��LU��sln�!c�8��Rˏ�	J�&e�	�qPw#6n�#�A��jk�<j��(�06 ��iwI�3Fl�S����{�����2��շ��.> O*�1����mU�8<��)Df���a���R�!��Fr<�*d�i0Є~
_�n����c1��l%�i�����J��e&mh��Bu�+��Z4C&�H�H�;N[6Lj�t���|C��k�(��pC޿6�jld���B?�Pg��N�6��q��}��c+Y����]�[Ȓ<ӫK}\�gˇ`��8�������	~�y�Ԏ��5n��aה��!��(u�����>aM�E�E6��S[�E���������v���e�E0�D}�}��f��&���ȹf� �W7D&Ga=�~����kq��7)�ۺe�"-'L�.{��f�F@i��:h���k�}��L���ݣ�f�Щ/��i~��̬�� s,?|�e+>�C0oTf��_��C.���<�x�5O���N�j��#��������Nd�S D��?)A)��^�DIX)6��ia}Fn����̘땉�KT��Dx��& ��wa8�:�=��g�rVm ���Nt�è<�孄Qk ��`;=�_��/>˰NU�������_�*d��YMգ�|!�;VLjj���b~'��.5�g��審�s˟HX)����#���
gz/l[JtHR�s����B���e���j`Q9�Ȕ��İ��V��n��FKY��kj�v���:T,� �����ޭ��ʦ�(G�����mY%���q,lkaؓ=k�n|M���N�����,ј�S6�U���ѷ�3��t��D�[�ʸ0�"3�l4�knr�u�!��Ok�������\�D�/�2cGf�,S����}���Fu]���{c�H'���ˠLj<L.q���S��K�G�k�0�A�7p+��sT�M�������\�_��(��tv[vWO�~�'9��@e
��
���rhU�_�����H�cMp\-Gۥ�/�2�^B|��O��9|��>���q@
�*~R�[�o�T�!�-ydJ�x�U�L��׃�}Ln�]ɯu��	ٽuD/��C֡ -X�a��	r|Cџ~[��[t$h'�S������3�̃eb�A�����qx	mw6���k
�z�l��^���M#̣E�uja����o�tKJ�H��r�K|a�#\���%����E+L�p,�,�+Ze��m��	)��s��U=UE�7(�_�2���s�ovJ��fL�M�$p�tt�;j��2M�鎯��]X�e]rl�li��Ne;)�f���5��8��T���%^���մCi<�]�t�nV6O��aD�
�����i+�Jru;O�Z���v]�c�6�� �$���U��u R�P����L^����hԹ_M�)�OTX\a���:nh�bao� ه�[E�5䅹vR�黃�*��O]Cs-T���7��̣a:�P�hf/�0����R���ոei�@�.4��[׼2�Nm����0v�U��M�N�G���I.~��A˪U���]@�R,�'�[Z>rtВ"����7��7Xm�D�?��zG9t��G���eұm��5 0��d�n-H�V�["��+ 0�:J{c���&�0u�s���h�l�$���r�N>�E��YF	���-٩�q���(��ω��K��D���f�c����S��Q��i�vj2m�M]J�!��� *��R�v�m�"��Md�&�����'Is��=���@��4N��E<I��'��v���"汕s[���������ff߄�aUok[x���~t%�>>p�5�Y��	�|& ��ӏ��~�V�T�4��ƔB{:}�F��=�@�fx�H�0"��;ll�T�b=W��1�9�㯤��щ��pL;dn�uA�
"�$�߼
~����O�P�4�tG��F�]#v:K4��`-��@f�ALP�+�u3B�T���rE��^�pa1�$�U;��ԭ������kwG���l�9���M�����$sC �O���ʡC�����x���p�!:�����TO2��1���Q�z^L�9�a!��nH�',ȡt������Z��G���}�oC�-���
~���;���p1G���e��A��=OS��X�E$.;�@U���0l���:�QE1�Zn�4q��"�d�s��-���i��?�� �)����ˏPB��:��q>��L[��b~�vڢ/Z-n@߉ϻS���bm1��#��	���]2]����G�AV=FmI���`�ߙ���k�]Yz��4#�w.��������K����L��Y���`����	�sA�L��# ����1P�{����U(�M�vR�!��*���%� �}#��ޞ�}3Yn�H� ��N y4��m3���b�!_�����{!1D@�6UՕ�,~�d�	�Ա{�	����;Y���]Vg9\'�L��HGX��H�ѶV"��;F�V�P���8"
%#畖�5JP��v��(ꡒs,F�'~�H��>��31�k��سzil�IY�*�fU�,UÙ�~�f��n�"�v�ն`�� n�$i�*ꌱ�Ȓ�����Զ��[OY���������.�	G+rVWV�����.K�e�����CC���a�� ��I &���}�"J�"���y�U��%�H��~�h�e�%ׯĤ��XM��C��p����ф������ۅ�i�5�܁�,_�d��%��H�֋ޕV>C�G�=ʻ�f4����v6�;�Oy..��x�-��}E��W�_�LC��B�X���]=�tZty�xR�S�Ӿ!~w��7�:U!M�4�z:B�|Ƀ����u�mꝵH��	�̓��O[�yM�B+�ywr��5�s�5a��@G ķ���4�Dw�&B��{R<��6l�4�;@��F��(u��������n�Í5�YKɔ�/C�
oH�.�{']Y��+x"c�/�L;�W��,�y�Y��	7Gks���#/u����¸k�QJc)��ۊ~���-׺LAEh�5�����c�Wr�yʫ�����hm����֭%AbL�o����#�;/>�VC��6	��#z�e��~u�(��(D���jvs�G{�� ]���I�0o"j������M|H~X�7�EV�W��Q�T�4�} z?ZF�SțvF���������έ�"a����g>�}hhv��R������1�VoO�-��w�̇��f�u{�Ca]x�%�u�]k2[��0��o�"׷��m���׃����e�"�S�	@������h�Iq�֬�7bؖ��M�Č�����ݡ�+)�E=�⣗�E���,�w�Cl�� fq��v�V�$�ʻ��w�Yj�V�`nb�啲�aj ��0�85�cS�<�
b�p��v��ׇbL��aq6�PZ��
A��i lB�$~C ��r��w��|��4;~��9�saH�-�t�\�f���7��R���λ�篒1��J����cF]�N��F|�އ�[��w���ɪ �u^P�kJ���y#yI�[�����k0�\�_d:i8�$\u`�q�uJ�Uh��xL�\���A?|�D�����T_EUggU:_{zV��+0k�.�#��7�~���K��d�FQRv54Y �{d�e�Yّ���QD9��d��"׾����k�v �hHX��E�	��Bi���~Y��_��(&����X�-��}JD�e{�Z�Ĭ)�Ce4eJzZ��ߑnj�B�Y9��'���+�]����L�Ɉ��Bf��g�����C}�eM�ɱDE��@wN=ۧ>�d�]�[
g�p��;�;�.��9D���h�WyB3�G\<�?K'U�R��Ù0�<08��x��͑��K)��r�tmu��_����Z�ƕ���*�G�s����B�Ĵx1=Ǳ�hG�֒>e����!���5�d�BB�A'�<i%6uf&�!�,��S�I�!��$��G��%G���P���uUXpZ] �,�u!xê�E��'23���Im�o�K���j5
R�'���D>o�s��ѿ�W�w�B�w�^`��+<�9�����1î�41�7ވjtKw�U;q����u�!WU�����G����pt�/�_��Җe-z�����ƺWbV4��^�n�z�1�g�d닇C�s�n�-p~X��){�^5mi�_��}_���$��Y����䮱q�p�+���4��^c �9��T<��c��xk� �H{����$En�b!����C��Z��L~/�vo,�{�"���(D:k�����cP������a$1�LCK���Y3�)�`(�_�}Ͷg���`o������L|M�Wg��i�i�#��/��,Q�����ߦ����*$��n���ib%d�Z�c����Ρ�ϰ�T��춣"yD1���kL�����n%���9�p��b�jD���-�{1��#Z	���`<D*Ȍ��C�f� ­r�<f�ޓ��f���Eb����]0�-ĽW�����*��HɅ���~��թ��yA�X���SY=Nk~����.�����BU�6�q�����;�̳,�uy_�CD�r�U�\��Y�˘��56��*=i�Qu4r��[���c�?��v���T��K����������` ���0�l�YqS�ؐv�F�^(/-�8V+�˺{�`��ec�04)�3�,��'-�U������n���s:V�z����>�OA���qy˖�Β]�Z�IX��d��j�#�LB�)�� {��"��zp�x���-aEvf%~���	�rɷO�E�@>��#0Bʷ�~�I�s���n�W�9�_���#3�VO��[6���h4���|�H���VoY@d�#�[	;C.��2���ʋ/z� Y\�1�lЈ���R� �r�VQa�Ⱥ��9�5���Ift�TcR!I���!2<@����p^�ҹ�I�.ŕ)(����%�,y�v�����N��
ߓ[��p���Y��6p�բ�O�%O4v\��P��Ai��{Y���Z��:@�?�k�,����:
vi������}���7β�	*YeVM����A���Iǜ��T	B��;_�3����3IXE����(_���ǩ�
(i�t�� SA�2�V�-Ŧ6	a�j�x`�*���Z�$��]veH�f<�k'0CpJ� �O�M�m#�XU�-��"���VFi���]Nt9 fv����]����͂͝}���*rL������~����=�It"ҭ-W���N
���6m/��[�}A�k"h���Zt�w�t�c�^]Nu[��z
0�^���{萿f5A�G`��ŧ���;o�>�E(kPm�Z��4��� B� ��P�5��4�͒2T���h.�Ŀ<��j�%�S��P]G�tF�>�R�I��x�H��{4֭9�S��)#��G�U�UyU���uM�O�����ř�7���[�R�<,�]�r�1]Ϡ8� 䃰�ٓk���p�� )�7=�k�qb9*m팃�-|fy<G:F�߻�\�����\��O-��Fwb:=q���j�3-��.���O�g)�������^��#�f�5��<��0����p���0�ﲕ?��t@C)���T�61ANk*^[���f+6�>���u���]�g�i5�7 �y��J��N��bƉО��X�V���:$� 	GV�"MA^��: <�P� A��}D;�����cR������0����`��p�QA�߀�e!ι	�ze�ͤB��7^eq_Sր�|��o�p���ڹ��VR�q����r��1�> Xr���(e�&V��*Z�.k����F��a��i����d�u?s�r�3�O8 ��"exҍr�c���	�!�S���;9E���:�LF���qmR�8z¿Ԩf1�8�ӊj���a!y5�%��s� f�J`�?hٍ"g����Y(��T� ��Br�"PP���~P��W�F5�:Α�G�?elz�Ý5�tfD���}'�5!��%+����+sPY�q� �_6������X�>$�d�~�"��>Q�7���?���r^�>9�$7V;0���N��,P��'��>ǹ��#*;h:�:]&J3�5���$5c�.�+�<�z�3>��i�����M�B1�$��"�J!�7+�t;C�h�1f����b�q6�1�jC��t�B^��#Fk����?�Mŀ��%�(,,'�e ��Be�/��`.&� �B����o!g�6���7�:u��l�NR��C�Ā~�*�cՎr��e+�x��b�7��X�u��n;ĉ���<w��T�48;�.u93.1�l$Zk<���J�Bd�y`D�����a�g#�3\�������-���ΝP	>�=�	��f��C "tO�?f�v��拴ǵ���K^��H��U��L.Q��-�.�I���q��ڸ��������	|��O.�2NU�����s�=��&/���%2,�����C_;����U���gm0#����l�״��П0ھ�?Y��o��H`ާ6L�r���J�&�f�Ւ��Ŗ��6��E� �#g�<j�,'�B��R3k�Nۺe��q(�WG)���j_W�ԣ�iOd�I�����)��@:D�9�v荫$p�ctΕ㶂D�y2��عs�.��I��u�����~B7d���X��O|�5=����в��X��JT_r��IE�K[e�
�a��w�L�Od��d!�ǜl�>��|tޝx�)#0���=��ڷ�m� eO�9ۇ$Õu���ŗ��"�����ū�g�#ea>8�F�:�>Q�4蚐���q2谐t���2[A�i&4���w~�:�|K���>��<��GLq_Y��?ǻZB�����X�=��&�R�Bkָv,�[�0�62���IU:.���L3D��]#�̛�D����[|4<EA_H�n��F��Bm���l��LKH���حe�1�s�������M�U1��^>��Ue$$PD3�O���k����O|������z�������_����$�P,4a4���{��~��{j�7JԽ2�|�g���cn�O�@������%݋#-�[�a`�7�g �xdNX�n�HB|���H
I �'�	���t_��k��T��Y�z��ZW��B=j�I��ф�\��b����P�e/a��]Q��cg��$��q����A��OꠄӥfW�|%�lm�G|T�>����r5����C��Ɋ�FO��y�QFoO/�f�N�V�3�¯��[-;}��̝��e-˙���Z$j7�m0�tC1_�?��`HD����7�5i������>TYI��j	�x H_���Q��|������M�w����Ȩ�^�g��/��[�N�^��_�Qqb/5��C�D�M+�l�dZ_�O�\Q|'�KS���g�=:?����}�[d�."%W1��9�u�à�Sm���V�Gz�J�9� ]�ms��g_�b9K��=ʯ@��u\x��|���1�\~�������;�꓇z��riv9�v�����s���կ@'�K�o�8��Ca,S�L��L�(�j~����5�O"�=I�uS04��괭�g�P�s-X��@Uɰ���g��0yh��~v�u�K𥿰�k�E�E	�{��4��`hY�����"to���C�@�4�q3�]��2u=�7h���N�<��>!GoF��T�EۇU�X9���zEIXuo�.a
)Ɣ���b�sF�=vv
��b~�!()K�ˬ���T,�D7���nm��Z+�^�����-�D��E�[Oln��c������:q� �Sx���,���fte�0E�g(๒Y�S�>k���L��To	^G������u�-v�̷�k�H=�E�G"e�@�5q+r=	4��g�/�\M�	��\>��Bw��Iq�W��QF6��t�L�3��Y.ȸ�n��A�{t���IS�F}��f�K�\`)�֘{�8d���S�f�B$�O��N>�Z_�y,����
!�$2���E`�OSW�y@�pe}8����w���Sq��͙���`��/��UE O�J���]1���R��+9LC�aB�ŦP�����/���tJ@��,�qd4@�mЪh������vI���e�3��;W�*g@��}�w�G�d	� &����S�J�BsPd*�����o%��r>�-��+��)]ә��cn�4V?�6/C��Ò�2��t�ȵ�x�]iz���'%����omC�G���{ڈ =  '�-y)�0�@g��E�3��[ut���&�ꈐl���	���DU*��.���#׹�3{�C�K}�Va���Z~]�z��J<���~�>�+J�\�'���t#^�_�qzj�pY K���Ip�?��a:�h F�I��f9���� �\�-Y���$�f�v�_��N��^�I!�[m�u:�J����~�Pǫ��3�άb�:K�2(�J�d��%k��eψ��6t)��fp�L�K�c�|)i��������,w�A�Q�|Tθv��0�#����V����skf�kx��cmw��Yz�|�� o;��E�������EG���GE(f�j�m��C�Y�~��ì���X�sd�X���5������g��J��=YmUDGs�0|zj�>��}`�Ms\j���jH;��͍�����1����d�J�Ѻ^����]��I
�-�r�+*L����c�(<�*Ӆk;��D��	h��wVT�������3&f��D�"cg>��:F5�ץ����
R�r(�WД��VdsI���Ú}���ԽvַoЮ�A��q��:�F9߻��n�'��K��{�e��	>/��JJ���p�y4{ e�BG-E��)JY˽A�g��J�A��}ŗ#㹐fj��-s�=r���l"�8��)��Լߔ7�9υ���[��9�/���6�J�������>,�+[�$yT����܄	��{�
cm��c��U����X�1[���Y)?6�A�M��^�
 .����1v����잯'�!
���g$'�p���#�yb��ESE���A^��������w,֥2Z���D�n���Q�x�َ%�f��^��Q9}Ƌ/,ԛ�6	��:�co�p��V�������atڄ+�Ĩ���#��w�׊��}�R�[�(����v�(F��y��"}զT�kC�]����N��^zgv�u��v������{s@�S��ooc���S$F����p���W�B+Ji`t��6?�-)T�E^��+�lx�M�*�����+��;���2&��(�Wŭ��Y�:�	���PYg8P�vV��P��ʆ��H�g�WN��4'm2�b��#7;='��ح��i��1��]`;��>u�}j��{r�K ��ۀЭd=�c�`����e�B�&"��Dk	����۷[k��v�q�໡ ]6�>?�Uf����+�*N,�΀�%��b]PQ��Qa�1��&emX�u��8R$�h�U�q�TY�Z�=Ys}8��&��lyMߞ�3;a�f�|#�y��ȿO��)�`�1�*)0�e�{�+�O�x��=>7T�{]X���x��Dt��0(����'"rZ�4M�K�?�摘�2Q	0��5,p���9(��+�]=?�<������d9��D��_�߫_�A6�<M`ȅ��Q.y�FR*~�	"	�y oŉ���8�����ZG�*8|Ic�:q�R�b��݃R"����7�jE��#x���e���R���������軑O��A�D!�JS�J��cز��m���(b��''v�h�#�kD�K���@�����;�w�3O�:��p�BT�cq2�la��]@�����i�ؐs꣭�h�w䊬��;�t$�a��C�ny���`�Qd7�	�^��ң�1�ݬ&o8&�t���G8P99���u;�y8M��u�Xe��'_����ϟF��	���;.�����cP��}��m��Rz��|���ko�0(e�m����5w��T���r�r��ڰ�
AG�������8�4B}���;��/�.>A o=W]*f���;x��T#���:�1� �EpԸy�$�=�N�eļ�;m��I�7�ę��l������ �LE,	Bx���/+-�01p�-����jpρ,��N��V���:�b���Xt�)'�j�?��_�����!N�/��8f���7~���,�H�hS�}�?`X��ꓲqs=U��)E��DV�$��E���D���`]�B���X�YO!��K@<)�3��W�� ��ž�sF��\C�p����1��Up�������T�	uɵ�iEm� (�b ������y�K�4�5<}��)p���{[eP��>��O���2��A�\;5˲�nj������{l�
��'���Kq\� (.�%���&�!@dW��`CQ�7d����Li�U*4�EDN<�$MU�ė�'RG����b݄o�^�r}�Ԁe�����������rcT;3�����GN�򎴖�)q�rޒ|��q]�xqЯ+��g�x���?*���<|�4���ڌJ�GS]f�ݼ�d����'�1�Z�YKI7+���2A^Iu-�E�a3�;N���wmT�^'�"ڨ�%gZQ�K4�Ͼг�M�l�(x��7˕�4��J�y�T0p������|��,�h09�@Ҩ�E�GP�)��z6�K���ު�����o��d+�L;�����d�ɺ^p��i[Q��%�`-���ӿwZ�k(�~�}�����N���r�����e�_ٵ8�^��t���ϫ�_��Cy�GS����1,�z���g�ƌ�M�Ią�o����k���cΖ�g�j���ɾ^r�������{Եoo-X�ڠݿ���9���Ty���9}:���6�bܯaɶ��P�}@N,{,��5X���RÄ�ؙ���W)�u0�,R8"s%!��O���Ȭ(��~Bd��2j|415�f�l��G#�[6UD
���Na���)#-�o��G��R�<L��4���]=�Z}����?8�>hj	���[�"��U�"��;<x��ew!F�0�<Y�l�V�*�韼-O\��;�W�_w���#�Vp������l�+�D.���H��z�)P���HOn0Uy
NP7��}�k8�8��c}<�T���L�����E�1@=��T><�愺��L�����~?�b���V��w� ��p.r�CV��(��Z<kF��^x�f�>,ݳ�*��W�"h�VBɛT��!%����;�L�z`��Ղ'(D ���Yx�,%�ŭ����JIɺ�@��[L�(M+-J�4�,M��v�ɡ}c9l�kH���w�����b�d^�'A�,���w�\(�B���`�/�
`�FPI���X�Q �@�'�}��!���H�5��~�>R_����t
p�>�zVcy3���Ϥ<:6�3m���/ PzCJ���x���x�08#(�d���橏����0�ص�g_1����4���u �a�Leg*V�Po�1��$S.�ހ
�r,ќ�2�7��es�ɷo+�A$2�M�Xv����垢��~|��	��j��ưf��E񰐅��~/��d�.(��$�p[������m�t����l|Ǎ�P&|la�J*[Nץι��{Y�f%�Y���!���Y%Ա��^�5�j����IB)mž��¶�����g'�:^(8vڃ��}�z�6��C'�AIoG���������5nU3����\6=q��zC�7�Kxc�h�]���ƾ_�=��7��b���^Dcp�ME���Q�2pV���&��v��R=���6��3��z�����l$v�~8G&�8T.��C2'�V'NGR�TF&�۞�Ou �f�?&"�9�}y�[�!��i]{���v��C��eL8U~=̈́x,�N�Ŏ�%:�Z���R+���h��2��7�ȱǙ
����f�lHX���v2�:�>�>8���Ig��v������hx4`ǅ�Jh����
[-��|�O��^��	�*^��t��j��0��� l% �?x<��E�V��y"���Q�B8E4n��+2����*.ג��|B������6F�_�y�{|~6J/��U3�H���)��@Ɉ&c����ܩ]������g]��Z퓮�cH�a�����6g�x����.����,��@�t�dC�B���lż��|K��]����
ЉV��OY�/� H�F�'xX����A2^~���-�7ՖX�T.۱ے	U�Ù�@��_�5ܥG�w�rX������%�NY�g��D�$�	�'�.�+W4V��|���(HM�nm*&+-5s��SjY���@1)I���\���/��{j�j��w��>Zq��Db���'�Ro�9*&����Ft��*�m�t#� S/ë��[t��eN�f�Ub��BE��)�j�Nx��bz�Ne~��LO[�O�Sh`s�K�ɂ�p��w�*�0�:bu�
�/�����q����.�F֫�Y�s��+���3k������F"��w�M��	�k^�?�Qr	Ǖ�Vp���u}�)Dn&i�FRHm#Ь��u���D�0�������R���j�~f���I���A�Q!�#^]vV�OK�V�� �XA���NAIb��ych�7X����&�G���D�;��%���&���-Q�ɏ�<ð����#7��܅�m����{3�~'�q�]GF�S�J�A4�{#�!��MH���+��M?���PU�.,�(J�K5��0�?����w;����"7=�Lol�cM�G�>��D�7Zs�!�)����6ݸ>���"��$����{p���`w���*c�[�l��yK�u"�a̤Y�7����%��X+�̈́�w�,��0RT�	8�D�F@��pg�@�W���e�Ǧ_.��蔒y��x�#�ä���A��Լ�fV�i,�X���r�ր0�.� x�0�����'&�F��8J��&c7�����B��`fqTUŜ�
7R$�&jq�l�ɻ�X݇�ŋ�� r����h�����Q�~�Z�R^%x��`9��9��"��<OK��|)��?�YW7?�P}�"(&ǬEFx(*��VZ1���t����x�a0<��0D�H���[�yܷ��m�}����ڶ����#	4�"�������5}k�ƬG�6-Y�o1���Jd��;����[IGr�A+��z�t��O�b���Kɟ��YH����~(~�z��O=`%y���P������g����f]5+�xj,���}�q�_OJ�/q����y�(�N	�Cb��MΣ�ͨa�D&03́aÒ�$���B{�s�X�u_���~:c��7$a[eI)�y���MuW�I��D�e�ӃQ`c��8�L;Ъ���\W'�:�������s1�|t2��ɘ�Y謪�
��::�vz�-���%$$1�h'M���/�6U����;&,0%�;�Y/:]C[�V�m��Ú�/32N����}@� �
B%�/\f���	�L1��љ�~�Nʓi�?��nm<~��#�4P)�"él[�n��&�y�a��45`��쥞�}��++e����+f_��J��§�x��0Q'ϕ(Z!��s���;\.�U�O8����/]���OB되t�cQ����/ރ)���1 k�%�p6z��<�;�Q:���r�d�4@�i�lZ]ݘ��Ǌ񎢿>:��QP���77��e7~_����F��y~�p.[̲P{C���*�����"ԇ��N�}�930���'��R�s� �l�]�f	ʚ�q���>�-�t���ʢ����9EE�ʣ%w�АXGHGfw8�l��y�<P���jU˰KsW{�*nS�� ��+��k��HVh����}Ez�M`��>�W�Η%0��"���c��xk�-��)�ru����,��kYX��px$�N\C�T�@N�HYaJO�,� (K����w X�߸������OH
:�%��Z9{�p60�)�/t�N������c��((��ι�rU�i������&���x���jc�f)ׅ� �_�F��+Yc�ﲪn ����A�;+ݠ�S.F��Dy���O	�00�z���>5�I��p��@ܶDJ��-�4����|����9M~o%�i(Tz����N�w?_��4dz}o���w �D'�D:�_+�L/BZ��:x~w�.�.K�N�㠢�D^�������R��j�0ƙÀ�x�L�|����O�[�*�E���;/񤂮��p�w�ǇgBsub�&�,]��z�e�1�$ړ`۞E�*1c
��ly׉�:�LGQ�%�pR���i+D~���K�|�/�v�:���ǐ%�k��kJ����o�<'��~�����n��g{b3�#��v���K���}�@�V}���o4����E�%'��
N�C��A��ɼa�z�n�%&�A���\���1>Fhf-�]�+��H�_��l�|��K�<"�:�)g�a���^]Z�F;��`�oE� ��90�:�u������F�ɣ_-x�#�A��s�A��D&�k� T��h�0���81�9�-ɻQʹ��Y��,�hhf:��*_t��2������x��*s�0.벥��p��?��BgJtu�+���_WQS�"��5=r�ɯB�� +���M.��	��&#�p��"��>������0�A��ź&��P�|Anx1��:6���cz &#Y���u���O8���P�R�BB!6hS�-g��C2��������-�����<!d�xN��1*�t�oXɿ���A������<��AE���6n8�b[�.*blĒ��6���1p`-�v�2�
�ax�p!DW��eMl^r��\%���Jt��kX=!��|~��d������~
����>'o��닥��^��xD�u�� _�]�,�S����tG�tH�#���1E�>hvf��~��ޓ��W�9�Rֿ��rQ��r��'-".]}�HF� �Z�N�G����e�d��#_��i2�i���+8�������B��ٺ�@�Ɠ�\�;F��|V����-Z�������n<N{����j���0e�:�gTV�vy�L�t�8�E�����qUa� [��Da��'���J����4�=i{���f���Rܖ�$�<�t�J���MŁ��'2֧�d�جhR`_�-q�;mG'��kǀG8��V/Cd�����DV��P��f�"�퉇�g9e�9�GMw���i[]�x'�u�����d�D�Ɵ�=�(L���d�{!�S()yl�G�	��nA�����$
�݊餐p��w���Q�z�����H(zG��:���^�e���
�O/oW�?��ڸ��>�����_tK�W�!y���F�0�^���snBsz����_�g4��匉�	�^�y�9FW�-�9��o�!a����|�M�㫩�m�pL�f�L�=i�6Sh[1E�(�:	���&�负B��~�aF��u���]I? �\1$�7cFw��g�bj	�x�,O�Z;p�<6��9��Υ��	�l��\%�W�*�UhU�2x�g��)!؊�&�5t�U3XK��M8���r�VL?Ŵ��À�����d �Ҵ�E��L�2u[P�ʊ��ކE�i<�!ξՊ�����yh�;��<���iڪ'PĄ�N?{�4KI�=����%-�:,W��|��ߍ��:���\���j7(@̈��A�(���i�z
鑽��g����P0�����=bր;-&@ζԤ�]��y��t�Jꛬ�=qn�I���,����֯+q�~"�{��q̌�qY�Hlf�t��qy��	��-4~���@�����&������*CV�Q������ڢ�Uu�a�<�E=/�o�M��1,�J��B�s&��Gܽ����y��7�ccO��նC�
t��9y�)I�5R����������:�MrZ��]��7Tu��j<�F�~ڐH��p��W�<��ǧH������v{`�5���T����Z)%X[G7���=�����=�{�U��+J��a�(6^��1�ϧ\�D9_��>.}��:8��#�� �.3I��j����ѱ�ԃ�|pqG�#���S���'hIۄl;��D�o�-y�6v�Oc�	��nf�N��G�`BFyM�@��vv(j����o\# ���A�E�=(��N�v^_�cH8��w��U��#�U�����y��#G���B�rV�`t(_�����dshT�x(�Q-3Y3��ڊ�=��tC��b�������\���­���*+�WjGۻ%�����ǖ��	�{clu�,�d��ܬ���M�lU�/ U�!��X��n��@��oCķT��[�i��X��@Oj��Xs��D�rU� R���xێ҈[*���;�	�>u�ü6ޤ�;Z�M!4K��V��o�'���1�!��Mc���U酓E���M#�h`1�X˧�e�C�������j	i0QՓǴQa���&�jO�Y�a���{��#>9�6�Խ\���r���ɸ��'%��F��E��u֖��⠆=�	
��^W�]6g��ڧ_S��_(ԭ��iO�I"����m�G����Q���~��iI�͵-�_6�"o~���^^nlC�a	/��C��p�������ۋ�ޏ1c�I����zUNV,����:a_�ipë��gK���]��%Q���{�+�״��I`É�R���rܲ�N�����.]��^���!��|=��t��G�5�5{-�_g�ħ���{y{>�h�='�czi�-6'� l(����6G�$�]+L4�=U7s�j�u�ڂ�5���Mr��O�s��Yo��r_m/��j4�ƛ2��p�%���� X03>�ٌR�
�<'\������
~`|�'�F�}8I���zp8������v��ɻ3G���E���rF�[*�����C������C�)L��~�GK��qB�1�p�Gl��o�V������a���eQUX��r6�T���M��!v�D��g�*ӕ�/����QŸo{xO�U\,|:A�'W\��v��)��Ax��}.�c����ȩ�Epr�'��\������_=-���y�=�6��dG��f�#c�,Pe�̣m��Վ�:�)H}b�����D��j�<9�@��	��PϦ��=N��R��n���[�0�x���%�U�������{Σ�F�������_) �����؂�dx-o)���(�u���^�yȎ (��afW���i>����X�O�\3��|�Y3�m�X�5����-3����=�m
��#Վ��)��u�}���[����������.aT|Fox����!p�c]n?�Dj��]�\g�V�������5ߚ�c���׌�Ј���h�s�ly�$pMU�8���))ۀwR9����;�\�6y�9@,�ޠ�8oG�:^�?���UFqI��A7�S���A�ǁwX��KY��3Ҹ��ӄb�O�tP'�?L�"��]��}]�E�6��P�]�y=e?��x̓#��Wc�W��_R�����H��ĝ�?�ew:t�KC��f���ƒQ�5S�~1���4� ������qD��o�*Ʌ��$){�HֽsӼA^����m��Y�#�鹉!yj5u<�4racb���C�� �}�&{ن�G
v���_y��\���h*�����_oיx�2Lގv��X�jzV���������b4�;D[�%�˨��-��Gvw�H�jb�q��z�����/�ϗ�P aK���.���M[Q���j�>/������zSBְ�Z�ϴ��b^&�����i�ڱu�I�]N��_�� B���$�V>Yh7R'c�����5�m��7�k͎@�fڳM���������h_�#�FK�Vy,x����f^�Y���ii��DA�'$r����_�߀Ǣ1_(M�,6ڹi���B��֎�/�1�c�P$��`%�%�ۼ�AD��7" A�=�k��B�˒��y2��6��Z�TB;kp�Q	;5��ۍ��� �m�[���PC0�AE���h]LS7���н�[�_�l<=��qsd��� ʒN��ݻ^�<����:T��/Ve��d��Ki�<��M�G�����M����M��Fi�%��E�1�;�-���ɿ���u��/�,O�^����U�·W"�ݛI�������@߀(�eU�`-�'_�ȱQ��Vy������X�rm��L� `���k��W�奈%�^��FK��<�����CA�T v�D@zF��^ƚ��?�R�q���4D�q�� KG=�Z֐�1�O}-�3�=��˼@6�H�;�c�~1��CF�Uv�&;�i��֓���9�^���Cf����N����'R�;r���:y:���Ɔ�����3�>�������Z�ĠA��	W��V)�>f�{�y8��L{N떉�a	��q�r�B�����F9m�-�
8��E������+��o��˸i-���|>�je�r�� 2�����c��6����%�ɣ-�u9R���)�06K�|�)))�=��"���q��>ڭ�b�@���o#�gr5�"��a��HM�n��Xfw��a9�k4�y��K�@�%W�}	�r���i��I�'ߎ/��%�*� ����m�Ѝ3��*]d��qB�Y��E�Ne��Dj��/=���(Ӎ��nI�v��,԰`'��{��/ ��<���u�%���9t�	�+���)[��.5�>�P�6�A|�LzG�-\0,w�"&e��X#'���隕��K���^XcDG�X�/$��?����up��[�^r��ԻC��Uo���i<�������7���-�rw�{��������e�����[�s_�4�9�A3i����x��Q�(e�^�������{�屮�^jEk���������9�I?�\��Pm̸ �5�F��O�I	α?E�2 @j]v6�2���ȹ_��򦘩��:��c��[M��uo�vn���!�<�4A���?c���(
��٫���=��̸����:��̐��X�8��M�夗%�F ��U���'Ƀreؽ��G�(��&�}�ֿ���zB��_vRC�8�\�G��#�L��W]w��h���Պ%���Kk!�x���hC���~��� ��w��kƏ�T,�(B�ɫ�Y���T�҄�`�e{7����
�;��&o�$�n֌�S5} \l��I���QvuQA�Ll_t�6�߂�V�]0N4�}�/�Mь��>�e.����<!�P���x䍠��:�]�Fܵ}_LC^y)o�&u��hصfaC49�k{XW���=��$&`����Ʀ�����S�oh����|4�ꉼ6Umc+v~�K;��T��
h��Y��v�����B/��y$�h�_hQA��ra������W~c��`=�����Q{����I�I�73��t@tNݞu�`n;�_C|�iۄA��B����yS�m�wRC�-����d�wҏ>�׳��+�}`ζk�ͤ���ܯ�S��T: [�;�'�t�w'l���55(�="�[Q;f��� ��/e�Mł 4H���R�;:'��¡�'����#�.������8�([~���MH=�-tȝ�W����ηX���͛� fgP�?Si�9<%.uYB��,�!p<FˌE��y��,FG��h�O�����KXH>I�e��i�`�{�3c��x/��E@s�b��Z��
K��!+�Ri B	t6��u5�;]�Φ���f�Y� ]K!%~ƞ('TUU�iL��
�*V�D	ﾾq�H�C ���޳�F��0�4�T%ݓl�E[�-f��H���d��_�:���ݢ��[�.����r���|o{���e�48�|h���2ЦS����5����Sݩ��g�A�*�����I���N�S�u��Ez��:��	m�Z���/b���B�M���4�hpUH�_t�!'\��;[Oٮ`����u��s�M3+,F3��}5_%"�=@t�\;RX��侷��z���H�O���P�q��7���s����E�@�BW2c5�"�TC���mH��_İ��E���>�Q��ŷ�|����a��G ���2�n��N��\�ۋ�2�8u�QASl������cU�+T���S�����|6u'Zk���743!D�����5���^�X՝�D1㈪4��\ �lЧ�U! uڭlc��B��Av�UI��;�T���vEy��[Z]�
�g�H���U���.�u=z,��NvQ��a�I�؊.��|uL�몍��p��I�xk��j�n&�̰h����,r(�V#hψ��j�29ې�^|����.�ʏ"�(O%���i��0z1E��jy�?�&o��`��g��0���&'��Lc:\��@���sL9>�d�n��Bw�ߩ#ۂ|m�+��=ѧ����Ը51iь�l4*!�d7A�������ʼ*�-Ԍ6�[i�h/���Ȁ�����R�%��{�jO��z�vB��w�m�Q;�R�#e���K]alτ������Dș�_�,��4�:���<W�J�?����L�r���[���4b+
!��W!�q�.C�ixXn����`E�O֋�B�_3(t���pr���}�O��+l��t��1z�t���Y�g�]~�_?�p;8
�n��0�5��4���򲊗�Ϋ��>\Y�(Y�����z�W��9L�����w�#�鸂�-k&j�3V ר=�q�T�y=��bG�C,�&�޴W%;p��^��GM���T_K� 	v�)�ed�n�!�t�ƪ;N6;v�{��c��@�ްSɷ�!�\����VB�E	� �'"7�O8�������
�g�q�f���^c��1��G�C k�٢�ř��1�"^�#�y�������%ݱ��xNW��]}ĵ4E$�"(�N8�y�h��@K�\�*wl�0Dj�`X�B�/��p������j�#����Ф��'��� ��
3��ͽ���F��踈W���v�H�~��9N$?2@�d�9���D���{�\�|g\��VT�A%Ղ�&XBi��6�E��cS�P|��]��j�s�qU-��q�"�h�W�Er�5��f��>�c�G��$X�8�YNoޒ���"���x{\�0^e�!�#4��qT���lzG���w�ڄ�	BK�OH��a��(LA���Q���ඹ��fC���D�z5�o��~��{��C���MU+ �
R��f�V�Vp�H�gbo-`�^�����*�-Ҿ�)9�:5����I`3��t��;	F��QC[���sv���l{��f�ɢ���PuZ:➵jα
_�a�y�@��1Қ�����w乔�p/+��/`|����q �a1����/�F􃫹��5�~-lW˻%I�Q��I94����*�BBl����\��.�9:�j:����U�c�)�k�"�4/��L iy��繠]��\O���z� fc��Q��M;�RB�Ĉ�s��cu.v�0�����2?�P=Q|�3"�2x�2ρ�/dת���*���h�5���r��5lMo̔ ������`�c����;��� :̣��O4�R'�+�=Vǟ:v�L��ɲ8p[M ���ޝ��ca�M�a	��ܳx��Rp����tMGV���U0�c>�\A|��pH�������#�k��R��w�/X����OD,rq�u�<IT�ӎ�אz�!�J~!�٣D��l)�j�5�A�B_�C��W�c�,�rc�d���ueo�"��C�(L�5��p�8m 췤�1��'��ز2��T��=1ܛv����S�{f:4���<k��)&S�O�vI&�z�@�Sj̛�����C ��a���"� ��:Y�*|�����	/�����O-��M����'=�%�dч�"En)�+�od���$�*|X�l����NL�:p��S�ߠ���Lp�f�^�j�5�i䏱�5���)�Ԑl�ƌ8R��A���E?ύ��(�1��C��~od��wO�@
��l3q��d��f�mzk݈z�m�FX��/��?�>֧�LD��?ֹ��[�+WL�BO�$b ���![�<�<Z@/�0Fq� K�;z"���\7�!�=p}(z�����j��$���=;-� �L@���ixh��G��d�njh�[˜��
:ʲ��x�O��-;Ͻ3���a��=,��������hdS�����4�LO��}���V�����x���j�����gz���K��(�9�o�ړ�Ak>}����F$X��P��B������1���%B&��W$;r?��N�� ��<Ko��W_�M̶]*�V?��Fƶ(���8�<2
V,�)�K�*3,�"����"���j�;��V��Z?_���Q0!n=�G�|�)0
'î�f�A#V���>�h��-�:�2fc�Y���ő��{n8����N|<`�J�X��H�6��7VRs�_~��WjE�����I�.���3���g6eY�|�M]�>u:-Ip0aä<�<�'��d�?���N�x$wz�����!J{���6|ۧT
\�_�&�c�P��Z$.Ф:
�w�\���w�G̣ X��~���8u;��Ll�L��]t�E�E�Tjh���i.����2�B`G��Ix�%Q2J�t�ܳ.��G=�A��:kyWO*ם~��}��*^q��F�f�n�Li��~�
���������K|�W����h%=m�*�P%[~d������,��&��	�#A��\�9��gB�Ik�5�������A9�1�h缨D�=#�Z��<����Nf-��%����4�.�J�����#�Y�N�H�Z���"j��w��a���7�d��W�mm�D(�pY@����D�OK�͖ar�h�w�5�_�&�?*��J����̴���Y���&� 5�r�(� �C��7�˵�QjIYwќ���Ep��,b���A�� _e�K{�>L��X�����9B��[g��	��B�Vh���=�d8�����⁼-;������$�����X}O;Z���,I�x�%E�����Mu�b��A�Ѵ��� ��?0*(�G2ޞ����!��c���0����n�q���5���=��U��lI��� �W�̖7�h�� �t�]�w%\Iƪ+��޽~��;x5o��A�ND�=y,,�yG���X��#z��3H.�����Bݬ~7��T��}M�-kPW�ot��*<�� �+L�~��۵|wn	9�0�::�W��l#iՖV��03���V�p��gA�vd܈89��o�.'a�4D���J��P�~��}&)�Uo��bp�p��,��;���~e�vȥ6	G��������(=RKd����{�g�
ܳPނaQ��5&n�m�����G89�G3�Pק-P$� ��ރA��5ۨ��@��B��D���֤�ޥ�"(������w�����6�]`T�h�k��Ը�!�`�Ů�Z-lS/�Q�P�����5�w��.*`��Ke{lkT�zx��q/~�4���a���y�a�ilE�bfG'`�Ѭg��n�� ǁlVU5U;�;�=
�E���Զ�Sv��A:�#,�ŕ��p�F�/�t�[ �9��6�����>_/47r�e܅�G}��!��E0�$Т��{L(h1����RxJS�Ɍ�!嶡�Z\Ճ�̍�!BT�w=l�z>+)�*]�{w׌c��_���Y��oIM`�}v�A��mY�wƹ0���nԏ�[kz���Vp>�=b�������ۈ�Y<�z�OTP��J�{DDg����C�4�`^'X(aZ8F9��.L�N|&	e�Q�u���oGقY����A8�c���?�cv����R�H�_GFo�S]B�ڼ)���؄پ̿���|<ϸ`��X����5h�@>UhA5�8�����pi:"0K�Oщ��h�1}��"�῏<��"t�ϩ��%��eQ����/���<Y�VR�*��u����B�fu�J}����<@��#ԭ�G�L�1R��6��j�d�4Kw޳��sޠ�~3�,aIK�\�w6h�6��WN�}z[�h����0ʬ3g��D#PR2�t���{��1VNLJ?�\�vcȏB}��֦	W]}����>S�A!5N���CG�:����HE��R����d��%?{8I��2�u���*(}aL�=�{��;�j�Et�n�9��Z�S�r��b�0���W�3N� �<�;���X�����wt�;~��P<��H���RS[�_qgp�*�����������c�d�4�aZB�����h<�P���i`����'&O�Aҕ��犑��
[U=�(�+��E��8�`�I���l�4���"X�[�8��άVB5��Yr�l+4nU},X����E	R1H�LK�;��{��!�H�o�����W���G��5�s[ �8���ٌ�(C�?>���� >Wm�<�X�+���'�V/!�3�ˁ�)"����l@~4�t��8jX�6�Ӥz�"ڥ�z� �Y설JW�����L��ū�h �K��}�pm~f_6苃�+%._�Ns2.�Y:��wH��ɹ-UD6N��A�o�N�j[�����X�ʩK@��yz�d��p�(�y3I)��`h�Gu���>��6З��-��&k `���_&�8�Lw���#�g��D;	���Y����|����o���ir{��ߺ�}�Ǽ�K1�$���qy���TC66��e��#�*]���M���qX��!�U�� I���F�6��5�8B�a��'dW&Qhº��ڐ#�<�����L�U��������R�ܤ���?a}y!�m���Jn�������������_:�R�V�׍���<�L[#_���@;�K2���6
�~]��)q(�6���^R�xv�v�[���e��e4�<Ch:)� ����n��]����դ�����D���hi����yC��D��X�@=.���w��Q���,�͈ݦ��h����ۡ�\�NB:���q�b9�0�)*>�����C~VB؄��g�h����չ�1�e��
k*·#�C��)���4I�j3$�f�զ�<Se|��r1��Ù)P��{W����A ��k�y̉V�7\�L��p��	S$��9R}Ƒq��н�rXX�� 	�
��~uI+z�z�:�6�_��i�1"S';�|$7~$&����o��"�
�O�j)G7��/'�������p��n5���A�G��2PU�Ѱ�"�3`꿓Vo��hG��ѭS6Lm@�u��@����h��u[�Oq���1���X�������!RA�jܯ uG	��D�gO������]a��[���\�P�WK�
����0w�^�Xz�9�č�S�J�����'S��u���i��ʓ��������o��]�fu�a�hO���o�v�D���%�n�n.�V9Lx�,gjn"��?��e���0�tF�ڲD?=�\��b}�D�kO6�a�m^�w�]�.�d�oi@��  �UT��ʷ^�v�y�ԩ�m@cV�$�T/��3�޻ �vQ�!P�mq��*���&8r�N��H�_6~��s��u�إ�ڨ�䤩n�T^����ի�/�s#����Ɂ�d���I�ׁ싴�3+D`ף��� ��K!2	�ɫb���"Ƌ�;�Ey��e�G���֞���ePM�S7q�3_Á����͸6�����߫�S"���Ir,�hZ�n�P+�7Dͳ:z���a'�\��|���3�4fj5�g�ҫ41�lMĶ��!����rKXZ�:�EB�����G��z�&����n)a�aP�Ѓ��N�O!����ޔء�5�r�k�"���b�X�)H�.kJ��n�!.��_2[�S�W��x�Q&���%�0)a�f�m;ɴδ��t�ܭ�	jnнn�?��$��-1��Q�L���V�.���:5\1�|E��6��"r5������by�pg6�S��s�_C�~R���`#�"ê25� ��\��[��֫M��s�O���u�� �E��t]M��>�5����
C���S?��,�D|=�
�� ��pC��l�A5�^\�p0ۣ��;���h�~ t�He���b��5_MڊA�`q3`�5�� �~� �/rw��eZ�����^��/}A�P��KpT��'��N�5$��T��^�Q�cph��҉B�Yo>'��@���jΕ��T�#z!����ێ��K���uv	�矈v������gꕽ�<mo�
�'zEF ?9t_Bn7l��a�"�%�*�܅��/(�T�'YB���|�T���e3��l+%-�-ؓ�mO}هMϾQK�XfY�hh^����+-{P{n��=�=���f���#P6l��FN��\�LI3b���d,q�a=�Y9��3!&�A/���L�+WA�%�Ѿ �`��c��Ȳ��W�$r=�6Í��}L�q*���p	s֣��Kdd�q���	��H���g1B6�3L��C!1�S���;��񆋧Y�l*�[}���mcϭ�ա���I��uH N��#���.�:�	�M�)�q%��&V�C:;Dp�U�(G#��\�-v
l�ә�{3��}�s2��ky�<�u�=���L����#� �9u�5�:�ۢ��goҁQ'��yE!��	nij��+u�py 2
�"G
#卲m;X3P��������ŭ�j���n��+��'����lV��&��u�~�{�Y�4��5|�6]�kh
���6��!G
9kf�~.�o�w�%_	5�N�za� 7����Mҙ��`�;N����u���u�*���i���<�����`!�%&\!�>�E�]�VX=�ϽSE������NBk������Gw��F�)��s ���v	$Ȉ<�h%�zW�����Z"J�!��tsV��ML�f�
�묗��iw�*��h�?_ ����o��F2M�Yݯ�4u��ݘ��gF�~\�jY�W>��J=�]� nM��j/�l� �����P���>-�������{�lizCRZ��Gx����'�?N3W.��k���4�<I��YpƐ�������C#!�<tE��'iJKa������Z@P��p����iB�zh?� j=���.yA r���dG�^��uEΑ:A@Sd�i�X����~����C��>
Y�7�j��}>TQ=ڛW��w,��(��J�͒��?\lIe+�+��N��Q��\��4�S��\��D�qdk������W}-�$@�uUe�I�c䈈
���2J��B:̏���q�Z~"g��� ��-v{�����q�J�~�(ќ��E�,�)g�n�V*Ioi^Z����0�UQsq�M66���m��jq
���mc-����1($wV���Q�>���ʍjM0�zҗ�rv#�u�{ARKƫ�/��a��}�(YG�Vx�Ovܡ�&	1W��<+a�&ҐOy���	�p���I��sE7�CQ_�N/џ�6���Q��Z!v��y�p�шŕ��w�@��6�m�RxVJ~4~��ў<ͼ�ؓ�^�N�P�<���_���rڱ����U��o-"�g$U(C��|6�~m�!M�v���p~5�n$�]N���S��1�9.zv����Ӯ�;��&X��1�vF,c�m�݊�R�����!,j�eB��U���,�4@��|J�~q��UN7�Cھ2��M�P����J�e]+[=��@@�̚}�@�Kn�+��mC�X�<t������W�R4+�w'��ТK����E���sQ�/=� 4���~�P�����M�� �o5����i�M�ۼV�����t7-�K�ޱ��F�})A!��yo�H�!�e�o)c��og��v{��g�5�|wg����B�G�}��w�o���V�C3� 	�6IC�>rF8ZNh'��p��)|���Q;�\]��k����wc �pvܞC������2�8��ᄘ`aS�E�<�����fRatI�>XQ��A���oN���ҷnW�A!���w����d���+(@�s�f���)���֧~VD:����_v���e��͉y�M�/s��2���rSr�SiD��Ѵ������,���`�1�`5�1jè�AI�z�F��ʃ���*>
P?{鯀;1�R �^eS��Z\$'�T���e�w��▏���x"�����j��Xn�}}�ߨX����
�?[��g���"�6|j�Æw��o��uT��7���|�p�lJ'c1z���M��^��^V�	�d~p�i5��:�oVNU�lyl��xb���A<@6��Q�z~=T�QC��=xq��5�� e;-j�
�0T�����Te���\��2�g���>���Ã���*��Xp�������Ri�tV��#`O��AH�Iܔ��X�&�-�|G�IL�� �n��$x]���Z"��!.|!��r�j�-ƍ�:��Ks�.4�c�s�
Cj�#V�ƏC]�y���t\��V<��H�5�1R?�b�e�uG!"(��� ��2��\�0d��+sY�>�'�t\ro��S��kY0�˫���<��ӈ���������`��RJ����,���F�2�7�{����{^x���<�a۫t50���J��iU2�|�4�m**��Z_�?�1����"�X���R�[yql�Ųz�21 �н�jy��E�Ү
��æ�T���)�*{P�5AѫD3��"r!+
��ЛvL�*�k���8�ě���r9�������{���6��b�r����(O� �F���&PLL)�gv��i|�⬬���u�Nm�ESN
����`s訂jȳަPpȳ��Ż����4�gH�baL������ƅK5}��(b�ّp��<9Y�5v�N�Q�ק�&G'�Yo
���ӎ��,i�����Ueqnl��ҨC�^���N0%�)��>~�����5�ڙ0����1�h�)���f�ul�Ͷ�&S([.z�A$��:�"����<!zT[~R������ECg�`��;2�{��_+�  N�K��Rż�g�a*ڱ���~%*�?o�����ٻfl��~mCN�	�W�d�b�!}��'e��H蟇��̽+;c7HQ6�,��[��qf<0bR��GE(]\����"F�L6��P�.JA�1�^���y�r�/LJ �@9�-੪zNd�m�e�w��*��B�{ :Y6߿��q���R1E�/����z��~V|����^�Y>�h�\�K;Bd%���7+-��z��s�Gtޱڟ���>7�$�·�B򞁳�ت�/�hQÝ�h�OBܺ����W׽)�ƃ|)�©�d;��Ū���j_lӠ��-���%{�F�W+N�Y�����m`zȦ@ݍ!Q,@��29�ܙ�E�cp����f�,NI�U�)�i�]�I=�''�n�7��R�K�p��A�WI���!_\�;,��bU�J��@���C��$��c �/�+U�|:�i�8lɩ�:E�L�_z|6��S�M5
�v�ĳT��']}bT3��0*ge��p�H�E;Nit���UsM ,H/H]#�d���d��P��� ���y��[���26�J!��/#�QyFݼُ�rR��|���cV[����ʼ8�v��Ň��9h-\Ƞ���0W^�[�Tt�?ME���K�K/�>���u�'5�����ѥzR��̭��%�_��԰��Ǎ��]{7ɖ����埉�r8����I�������6�vY"Nc����֥ x8�	;�^g����崩�)��S����']+�>��Y+ѣ���IJ]�[��	�C:אָ�/Iu���Ԭ����8u��k�e߂sy苑��O�S�C�ɼ���BJ�6/�v�*|)ذx�)�ӕ�E�z�G���B[:�&����é����0��������e�T�r�)N�{s�jDj��[�F+s*��iDe�Zk8lx+�� P����4i��`�)ݪ[.�B?�H�흈��_+�⸏�M����� ���,T��(B�0��a(oѴ��֒���F�OmT��Fae��7ãs�����}3.��n�ɇ'�"A-wf���;��cN��~}��u��ݠ�,�k���*dyVf��J��y�&��A�G�z'�]�e>�!F������l�+A�N�B��iz>IT�s�˭��i�k�h��l`����k��|t�]�(�I˂��@���*Zi,;gp��a�nY��U�v}�O9U�/��'(@�Ȉ"���v�9�-�w�k*N��Q�T���RwO5��?��ߐh�,�,ʂM�Wi������(o���BZl]�&��'�
��b�O��(�A,�!/:�*��J����1�ӓ���ч˝�po*��b�����ѓ���ߡ#s���Ո�J��4����N#�f���:R��h�&jc�e&
4�[G\,���<iܲl;���䦽�����_gu^�Ƒ�zAɱ��k�Z3���Cs�ʘ��� �`��h�3[i��@�q�$�_kJMx<��}�ٙ���q��өp�@���N7D��H��-����D��Q�����g�{����P�I��qI�Ln[x#h����Ď�Rj���c�u��:
�{Ԑ���iA���UN��d*�'V��0 t�>�fh����'�bw@U|��;�]���L�;�9�M��>^�x�4UVH�8�glȑ�*9��M�X�����Y_<�N��<���=�
�̋%� �� ��[�in��yH�%$66�#��M�AL�kQE.�;?q�!��.��{.�$A`�I��4~jz=�2< �l�]�3D,��KyX ��VP]sW�o�F���p�6I�ŇT�`��u$aI]"8��)v�Q@H�T�I�M��߁��녊 ��c��IܣJ��(�o�(��S�Gk]O^�T��׆16@Z�-�9��f�iU�Ժ~�`~bz	=e��"�x�,�d�vK|RJQ��7�sJi>5s�APs��{oðZB����<��{B�����YxUn�^���d��#X������j��Y5���ŵ=]x���Ul�a۸v0ӫ�&� �fX�ۯ�{�c�l#�U=1CN�眸��"!��e�?4L�����N�R����o�;�j�]�F����A��"T.S,�Y4p����37��>�o�GFj�yw�B�>]�~u�,E�SO2�I�=�Or �~����H���-����uf���?��/�a��o0m"g*f0$�'��p۶ �z鹑��E�B�`�/��O���l�u'��<���y|�6!���O4�0���f\8�9�i�����몞��raW��8��i��n�7�iJ��� �2eO>W
��`�re$�x�j��'O�-�Ă�S���� ���\��VB�\{��ɋ����g{n�?��8:�6t
�ۃ~��P�o��*��.��0���4(��i! ��Ŀ �����j-ׄL\��lu�#�y_�_��c�@cr5��[����H��%�(}-i�������^`����)2��9�*/j���^�Y �#�A�e�I�C{�W x	:zV�)�<7 cZ���`�:��:b~<\fϿ9�Ua*�8��/ǘU"�0�����#��tKj��	vmǫW�՗F\�<�D�ʦI��=�Uֿ�G�.6��?���j53��n��H/U�S��pJe������	fD�uQ�f|y&(�D#6pFd��g�$ xĤtj��t���Ѳ�k2�{a}�{�Hi�洙_xe5����h�C,�����n�g:65�M���AHƬ���P��nT�h���y�E��S+��[���Fy����A��>j^XK�F�m��Eo�$�:��0��I��a��_�?B�Ce� 0�ۖ��_ʼ���#�"&A���Q�F}/k�����}O�=嬵N���S�  ^�u�>�D�Ďu��FL}���Y�.��^���np;��v�K>������3V�(��?�=m�N=8vF�Mm����Q<.�!-?��J�c�K�k[c����� �y�m�`���f,&��*���C��.���̟S�&��+�xz�C0�� C�`*ї6���v[)塐�`�c���B�R6�n��p�M�@�5	�+h��ߑj6$�'J�l�s)�x�Ķ����U��9BC0s'I����ĦUδL�Z���%�����k!Q�7��ۛ��JR��mE�(F�kM+\����16������.RmI��ǋ��P#P:�q�O�vS�Ɔ��M���%�11��AR��9����*��a۠��, ��@ �q�7	�E��E�v�+��.�2�|;H}��`��� ���1����*�*����9�F�� |��K%ʫ���߬�v|ʳ��Sm��׏[�,<M�u�º��]�^�5B�yc4?���X^ue�L� �z�d��bS��T�¡��%��?x�ȓQ̎mWE��k}P�,U�k���s!Q�b�S�1���[�$���f~�ҺQ�05�^�{�[����s�aIЎMx8�l��~��&�f����}W먀FC42��bj�F_w�I�<�wC�t�A�	]Gs��o������dB��}�W/6]r��l,%(~-dF��!�W�p�֧�����i�������<�H%yYm7��j0�V  ا}�L�#�ɏ�U��P�C�#���T+X�Ґn�Eȥ���a�Y��'�@ǏVj�N�J������nN��{4�$VbrbZ�m��L���p����J�� �0��_��zzQ���.l.��y��[��\:E���_G�8����/=��q��rMm�ן�$�DFb8"zW�h
���l�[�E�%�����K�����.̼��L��&c�Z�'�+��6�Et��?0�o�ߥ�@>�׬v4�2H{t{��0�@1�ɆS|�ŷ��D��~"�I�����X���͌)�݅�|VC�Z\q�=N��g��@��|!zڸ^66 �A��et���̼hfݴ8��,�/5�b2��.8b#����MF���Y4�,�'F|+�֎���܆Y�E'���խ0�+�*�#0����{�O�y�Y�&�١��׌�zۇ?.M�ٳ|	�h���N�����9�!�_ā��}��K�fҗ�m����XC�{���*P%XH������9F:Q�ӵW��A ���B�Ll�����er�[6(Bݸ=h�v	�̙��Xĳ��F��e&ٿe��7z��n�s/-����GA������q'�/��	� ��ϊ����.����ת2�-	:Ć����o���F�M/�@�6���
�Q�3C:h���y�"C��N��_<0F��:w��`s~��%ѕvr�9��~��A�Q�,;����$�`�9d�mnL �0xJ�@ɠڻq�}!�Ľ@�iI#��ݏZ�=+��X��/׺������yd�Lq���$��������!Q�[�i��A�쒐��'4�:8�����NL=����D��n�H�5ޅ�[��&G���!�T|6��*��{H�h��ͻ�W
��x��B%Ma�!�lq�W���"����l���䡶+�$��쩣����I�H�=�D}��i��Oێl��j�}<�5��A��$S��Q+Q���!�a h�x[q��8��p������v+'��1�4�4�dIg4��O=.�N]�t��㖔�~��d����<���� ��ĩQD�6�S<F؏@|�?nGz�{�:Ơ�ڱɔ3Yz�?Ô%4����.�����""P��4�P7L[�Og�`2�"��F.8{gљ�Q����T������M ��<���}�-�Yi�����gk#�I�&���r�
?��Μ?S�5�����y�gYJG��M͜�A��qX�/?�/�e�s^�����%�γ��4�c2`�0�瘢��������e	���a?�S)���\��Ʋ��/b"�G�5��0P`i���>��70��q\��=5Z��@x2�O�}��8�������'9Xc;׆��^#/I��Y��������z�b�,)�U���E_.s��&DN�G��O�VR0��I��j�n����`��&��_3\kwD7�"��U���L��`h�C��F����\�ζ.����e�,�*�k�X%���f�+Rai�U0<�
$�uYO�ļ���K�$�^s� ��k'�|�a<LR�H{��%I�Ʈmh��_�l??��o$��@1�N��|��u���혦%BA�������t!��L�׫q�����j*�d�P�-=���R��/��6�����<��]6�\ zQ�;<MN�����}:[����sxs�g��;�� &lvar?]��M4�|��鴟iŜ�j�Mͫ��Ia����YJ$�{��6<y�����Z&*D��<
��I�o���� ό�0N�I���7N�	�Skװgҽ�+�D톸�����B�*�DsI |o��A�"t�+��@��R�&�ݰ*�2(�Zj)_���qj��b�>�h�>(/�T�I�."UB/2:���:F�rI̯����O�����-N9�V�R�&�h�0���ŐT4�#�"�/�F�%(��}F�!P�@Ů����&��RD�׽�5o�$��(�ܳ������q_��&{R��ƥa$f��e�J؋�K�j��YL|�������҃�S��0��t�]8b��&��(l�i�liʅEuHW��Nb��Y�<.������b��%���p�{7cS_��f+�m��7x�kbx:�('v�	����h�^����z��<Gn���K��?/ޏ�T;��xs�.�I��@=���^�7�~��f
�eX���}�7*a���Y �l� k�[�>��W���c@\;6��u�B�����ەڰL�Q>y,i��bB?���3T���������9f�V�Zk�Ԁ��0����&�I�����6�6%��}����1'�L��"��������1X��3%��l7;�Q���y�'�t�������"9�7�#u�D�W��$`��[o�WD�V� �A�J�77/�Ių3]���B�y ��hfbt�wk0�O~I5���/\{W�P�P���a�kDC���Wfx9N�N3�M�tX$zzDY�;�Q�IF,xOׯ�u��w��ѹ�H7hP�&D�K����%�넵1˅�6�������X1!��3�(;傈�J��T�_��N��x�T�4	�>�V*�rҟy���Hn�ĳ.��iW3'S���|1>������z�leڈ��~�SԆt<�m� }4�$� �`z]EO���H��|oĶWu��G����g��������@�)�B�gt7V�qwbq�b��Bx�%����a���.;c:��<<T`�_H��u�p���;)S$,��SnHҁ�˰���������9��:��哈�_Fn�Q���V�'`ؾ���%��B�mO�eԱ�y����J�.G���,&��[F�+��$���ͷf=>��~��&L�d��aSy��"71Ü��)
�9��!*8���;�����y,�l��=�W
H=As h��C���5d��g��e�YEF�h�\�ھrJ��/$��5<g�8���(��|6�Gv�}e����=%d%�Z��H����&V�����,�ga����-�[��i�{=Z����_��BrYS
�qq��؁u7�2�J�����YoW���-�P)�`�l��V���.��C��)J+#��I��;��F83�C�O w�!���n�H��R�1s�|������L}Ky�F�a]�>f��N��:�!�d�>!�6�#N���r���y�A�x,�C�{�����I�QW%\����GG�����4dRqV�K������Μ K�x#��~ H��,W�r�0;2NK[۶��<��<��xY4��М4rs��}z���Zۢ�}@1u��#��Qf�yjl����Z��'��ael��	f��� ��h٫���	�\�ք�r�+��\?���?�b�cY�� ��xЎM�1�a�0�|٧�n��*�w_�dݰxv�f�@���V9���G7!�Sm(`�>c���"�A~w�8��q��ֹllTH�6�:gH����3J=k~�ʕ����UQ�5�a^[���?����u��R�E��d��e9�|��ּ�KɞP��M���[4�s�䩌��'jFwR��|XЦ~����0��ֆ��`��E�Cr��qd���g���`-��88sf��zi�W����D��}�+��>��Û��/��\��x�Q���O�^ҪP�I�h�_o�bhD��07�����O�_��|0u�}�_��6;l�a��e���x�$�۪�}�c7M�M�����ęd-.9�k���߄}%r����`@S��x�6l��t���@e�eG��m�P��x�u�Ȍt�%�U^2%�z;Q�^����V� �����;[����'�BU���|�u�ݐ���P ��f�'D�b5�p6�*ֲ�)�n��J�zpi��DM��]�z�7,��9߿pڠ4��O��7*�{_9���`�w埜H��a��\�I�5��J�m��V��i]�\=�zJ ��0_� f�T_��Y���+�1TXz�Y�6�qz�-Q}]���q��b`�Ag�ǳwR`6 �2�rz��@��B�|�������2�b��_#Li�vV�P��M���\#К����f1K�Q�;u*��/b��ͽ��ʽS��,�&h�˵�Ac�Mm�-n��g�g���0�魟S���3O_��b$�zh�o�`]�b��u����&�MP&���ׯ	¤/)������7xdXt|FO��栨T��6��k\:Sq����P	P�l�<�@��Ix�)���0��֘�M�`$��2��r��N�.��k��E��4�nN2�r+���Yٝ>3ѹ�O�r���x:�i����]�E�s���ҴdYR3����2V iq��'8?pVwۙ�M�T�j�Ù�Ǳ�P:�2��s)������֕�J�t��h��l���PƹfZP��=�}���U3��+���Q��i��P��.��`�ؠ�roEA]�0�)/�VեjB��G7�F�?��\bɉ�L�)埍������-�Ɲ}9�����2E�M��U�VɭJ�
���������g��
8���%�OL����J8�50��>i}���u�.0U�A�����k�@
s�<�
����v���/�Tp�d}�Q�`N�xEbT��K%����w��/�rxE7�Yр���,�D �ŀ(,�-� �էlK�xр�v��`_�@��&-���=%��n^R._�p��+$ga�z)ϗ7҉P��U5�EmwQ������q���*ʛ������A�@rG��㭠0�{����p:�'���7�����딞6�p��qt�~�cƆm���UܖcG@���̇��2�o$��5Ug�FQU.h!�qp,��I���/k���r"��x	��.�ɦ��Y wr7�� �ȗ���Z�r&v� �f�畈K�d,f��
��=Fxģq�߶��0�NYk�6Uh���"�YֹG��#vLcɔ�e@]����6���:�3�)�������-t���'��I!iXI�on�S�篟�I��Cƀk{���-�M[؃g�������M��u[��j�Ԕ�����5XZ{R�����EE�?�S�(JgU�oX��I�)�-J쌃m��r�+�K�&ה�v�k�@6*�cA��$sR^�`��z���8�
�"E��u.����r�t�j "87jX�{��G�W�
�0|9���4��-˷�G�s�^Teպ$�saC#������0�r��Iz;�?�Fτ�$�P̅i�)�O���TyC�c7ay�V�-G����\���lq��K�@p�!SrT��A��9*��s���g�F���h��9���:�ep;t�"w�ѳ1d_���Ž5ɕ��(�����
�4&���d5��/�*�o��꡷5�]x����D=D:@Bܔ�>��!�S�ۏ�ܻe8	:����}�*JdsC��pŭ�̬�XNH���+E��	Nk����r���a�Hh��y���߮~	<f��ŴQ�&t��T[5\z�R�N��M�$?-�-��/U�|��eB� ��!AA�VמeI ]�>�#q��f� Ch����k`� *��m�pV�S��-}�
0��#�{q>*�ډ��o���?t��UM/ �F.6c$��;��4�\�e�E�4���kA����X�+[(<�v"�71o��W�}	}Ȕ>|$����Q�����&&�HUPCu�cZy���R�R��1?G\
V���K�<�`@��zx�t}"yh��n%�u�3�&�|���Zl:��L+
5�/H�l�P��i�Y�y�!C5[m1�x�V��v�4��E��e,�ߓkT����7�t���-Te蒾�����J�F�����x��$�7A~X���`�iK3wՒ0�W-]�/m]U��+?�%5�(9b/���Gw�6����K��%�4���ƍ)}����l�o��Ҡ׀�bR��H_�T����^���I�r���l�/v�f-ܳ��8���8���9`�֤Lhm��֌�'{[�c�H�(�.rx��@���<e��o崮!�G�����c�b�l~���>ѻS���RIRE���'���o]���Fpq�ӣ@�� ��B&;OH^��#M���	29;�3�X!��u��Ti�alYx�^ʬ��Z���z�4fNΎ�G,�u��i��Gw�7=]J�ʛ� 1y��Y(����P"��Si��m��;��H�No�d���QD-j���<�^w4�!,�8�*F�	�&��'S#���-�jT|>ɰ�&������q�h|�	)����Җ*2nPR}�{����mo�hGV��;��!q�͈��k�}OrL�2��L�i�~�Z$k��s�PXӏ�	�:�$�gf���A3��7�b����{�?��� t�K	�B2L%"���8�mB~�۪)4�*�M5��C_4ڑdG�#��/�M��Zo$�dh8���v�"O�؊|�ͪ�,&�7Ԑ�-�l�e��ɣ#敩����D�G�I|�	��O��<���8��HHg��!J�R��{^���vx l��)��u%��s���.��5�ŀ�Ɉ��$�Κ��x��v��_�(��KJ�8��v$�d�����1E�ߞ���Q�������%�Nos%��F~�u����s�Rۀ�>�R�n�̪{y�_�;X������-���Ękj[nN(0��"�)S[M�ZW8B����Q�J��\�섿�іf:�h��ς��&>zo���h��b5�l�nS�~�E$�Yp7G+N8��a
p�U\꒘���s�＊aEAW�^��y�@?Qy1��4[ؽ�Y!�:�-P�ȷ�>��\���
J���#%���nB����U}y�&�"��l��|�t���'Č�F�ՙ��]2��wr�a�Ĳ���c�B:*��6���T�,�z<���歝H���!�`����x��|+��{��<?7�dX�8�M9��O�p��m͛�a����O��~:.���fR��#��&�x?A���~R�0׎�<�].�2%��f8���s/��H+?zY2�X��p]��?����' ���/���)eǩ��ο�_�OA���6�H�ʪx�/ÉY{���Dp"6����Hi:XaJ":���ɤ( �#�fʳ诟	c��k���_(�9��]}���
�y+�>��q {�/�<�tO�9OW&ecpV�\�~���b�n����,]#U����d���5���)�b
�l?����Cև�-�_yJ6,T��Y'
/�I��G�:�?�lӣ�!�F�~�6�������:����IC�����1v??MA�2׾��G2����M�a�Э���X��N����YE�@�A���GT��s�.ni�=�������ⷀ�,��U��$є�����Ǌ,�W�ό\����Ց�h[_K�Ο|A�)��{U(c
9l^�U��Q�h������V,Q������^q\LM����guߒ��iΦǙ�"&���{Sc�1��oGĝ<�c��2�m���j�A�T�q��}�xc����ZT��j�2o���i63���Ox��>#} '��f�Q���L!q%�݊��0so��擓�Ā�8/�� 
���XI��oxw��I��/���[���яZ�)����l�y��- ��"}��.
cH��q�m����r�g�f��M�{\+V����%82���+���������6�.v*v�t-�75[�.Ǡ���)�.]��l!>��2?�`M �7`*mI��9^��y�֙��Z�Ο��N�� ��dQ�0 ��Sk�S�&uy�:�Ȋ KYBt��їǅKd����w��B�0.���"��pS�/��h(�?eV�)*�%�Rђ��W��(�lK�oDj_� P���Ȼq��1�JP\w19O`�$d��k埆��b�Q&�v��캸�μ������-BH���Sy��)���P����`�ɍہ� v���Y��.�I�ϫ�5�U���5���jY0�o�{�v�.�G��Xг׹N�hQ�g��7�H�Q`
��y-a� +լ���xV�ub�*��FA
��m�em��T����(�]E�t��g��3`GB�׻��ˁ���e�C���ZH&�yF
B�W����9�4����Q7�i�:��Y�-W�Se�7q��"N%T+�<�P��X�U-��_:���p6���M!��_+�ل��Q#,�N:6ơ��T�vB� ���� O[ϿyxQ!C޵(���7�����+-B˛xT��[��[��h�0�&�o��?��	��$Iγ�j�O�%d���y\�1�o3���=8+
��6zk�Xs����{�f!���<�S��,2<f��2wkD��s�R�V�U���[�����&��I���˘�U�G�h�-�٣��Q:>����<&3?������L�ͮ�s� ��w�Q?/��8z�����Ѩ�\��W��^���	HSAAE�ο��=B'vt��J�1.J�S��򱬜z:�����}o�:��
��/��m�����H,5W��
h��:ѥ9�w,��G�G7��;){���	�G� UK����Q��b�5��6���_�̸��݋�Eӵ���9�h�1���x��?g�朅Q�˘���`ՎS�`���ZO[��^W�?7q�Ro��	�OS
B%𩑹U�	�G%vY���Z*c\�
�3��"T�Q�[������}�� E�NCi�����LBz��Zv7=����b��$%�R(�����k�����|���*��� ��b;`�|�ˇ�#f�3~�]&E��ȭ�����|ZL�;~�{+E.��^��#�҅/9��(F�B�z��݊�г�\��ux�>��vˇ%|r�Ȝ3ߔ�����T�mnI�wff}��~��N�+ܻ{��#��g]�O���j�6�ܘ�]c�����:R7}�8�4�@��&d��"�Ǘ#�X�v.VB��8(��Y��eG�cIm��܄}xIJ�;E�֖X�}�����p�d�ƚg7ף0� !+��vo[���TB�������i��։1Ȑ�$�rD?G~�4R�M��Ry��GZ�B�70r�N��7�i}��1�y������>o���� �V-�I��t\g�ݜ�/b�X��@if�B��W�7���<y*�LT�R��b������y]ÇK4�oL�Wan���k��{�+w��\^
�İ�P��lr��
���!��ԯ $�6	�$�
 ��T��䯫ҽ��\���%
�A�.N}&�v�SLԓ�~��>��	�[~a����}13,�Aɢ�O4��="*�QR~�_^T}�+a��<?��{�m=�Q�A���>��+�D���X��ӡ���Ѩh:wj��~2�<Vl#�u�]�����ן�+��@�Gv���ѐ��Y����Cv�7�$/��ql=G=�a#AK��
��������WG�'��)��<g�l�8RHx����9$�a�f�~CR+�C��X�s��6\wi�<�)��)�P
avjF��0ZD�5c_/	Rz��v�U�xŅ>yR�	����B,�����p|�2u�Ha�Ve���o�O��$�v5�����['���{���c>�jR��G���I��x�w���%�U��'�O�R�Q#"T���5T����@'V��;y�?@bT8�g��I����>�ۿ��&�K';6��,��୸���X1�1���8�L�4�E��������� ��Ot�c������	J���4�7������U�b��?:U��w�Q��u�mc�r��	��FJH���Ma�aP�lݱ����]AT�]��c�t��֔�a��I�o^�o�5QʦS@v��u�6o��u�qN_��R���;D�Vp��'\��]�w���C���r7�7����Q�tA-�_�(���!7�!�H�5)�|�e`h:ݪK��V.L��^�$���=[��%���Lv�Hw�9m,�ncu���1���t.U�b�RCIT���n�G��3��+�Ɏ�F�s�ՆO����%��!Eg���T����6xfb����d�ԯ*�%��e��K���H΋lu�Z'�"�hjp�z��_�&\���_2�#_1�zڡ��&���l*8Z�P	^kn��-�j�),9�u~��?�Vm'��N鿞&g��,z[��[c��e�w��qd2���d�2���싍�������
�z�#�V//>����XNj��a��+'� k��M���zgd8��7�n/DA`j��fYd�r|��z"wz}��'Í��P �������S�I�b΁��5󂬾֥K�->�?4�ն~�}to)W�>�\rcâ�� �1�j�>N*j#�.�P<��6�ڮ��1c-+o����N��W�ѯ�FqU)D�&�j��c���`��=ظ�6��T��0�G8,����.�7��^p�?4_<v�DdS{v˭C*4Ce�!���qss��l���2g ���Wr-pgP-�F��M$Z5a}����Mұ�����1��3n-���� �ˈ��,�o34v�i��)�B�{���ӴN�i �*P����#\y�=5o��Y�c����_:����OV��vޫ��WV�������#9bA�����l[-��[0���b���9�/��0%&��9��L����� �-��x�W�f��/��`az����f@��^��8�݈6%6�7��p�	��a��1S$��5�gWK�h.�4� ,/r�nݝ���.8�_���ԩ�M��47$��x�����J�/�괸�L'^>�F6��Y�d\nd ]�W�@����>��C$J��!���,�hF?D���[�U�r�&��}Ó���烏pN�Vì?��GO��Zeqb�'�VG�m�tc�ÔF ��=u
Fz�d�E�K�|:�|)�o����ob�F�5^��0i�;ߛֿ7�1\`��m*Q����Ӳ2��o���4�{�Y��sqϴ�֥/V��N�h�#a#
<K�*�R2���/��M�-«URS�~�kzk.�|���m��;u#���A�.�,s���n%_��:�7e��&@�H�=C����jb�K�|����[��2�v���en!h�+��h� �o�r0L�{`@�QíU�V(�u��
K���#pem�܀��#��"�*7���D�Ǭ��(��Z��G�0�-Pz+�f6V�͈�$����`��M����+�.e��)Ȳ�:�ns�6��G�I ��[i~�"�����
ͬ�n#���
]Q?�	�GL�/M�:��6�ߙt���`H���r��L��3�c\�6��_Ƹ�̚�u�̶<$�:"˥3�����C}!]Շw;�,��W7����^c��xPT�=�G�Z哴�d�v��E2�$�����ȓ�:��CH�zNţ�tE]6��������Y2���U"�чl�K,����3���ߙ�O/~Ҷ�"-8��{|J+�0��=F�ۈ�LH5�L�.����}̵K���d��߿1�\Q첮�����tD�����x��� �)�p�H���y�
[\ x��Ӫ>�b��5��LF
�u�����&r؍�ǔ�i"�w�n��1H$��)+�CV|��m�!(��/5��o�⠶�2u� �M�FvҘ*g�Y!��W aXU�
�[~,,6�l��cR�����8��+*7���+�m�ι�utP`�!KC�t�Nӈz�4<�A6?�	��B��I_���F�<V���\$yv	&�C���k��6�<���X��76�����;�taт��ܢ-�����u܇�r���JF�gǓ�&�wB��w�ũ�PN̲_A:�K�+�u�����t<�M��e�e���zۃ�L�y���{�X!˼>0��5_C��s���
�`��?F�y�3����,��������8��uL���ӷ�WZ3+閆�w��j]���J��pp����L��`��v�/�=�_�q��`F �=V�'�'���aMk�=�j�L���mnv�FE8���5���=�T��\�Ê����?�e-�28[��ߟ��F&��v��Kf(��Yt���&�`����Lq밟5������_n7���$�/���Я�=��
H�T��5{G�8择u �̓D�y�y����]'��sHTb��@����ڐ�#T)tV�y6��l�w,5	�i��aE���o�z�Д>1+XELރ6��&��A,;l����k�o�C���%�����-�&�_8hT�=���r��Ice�<���x3s�{2c�"`�K�G�^��,O�:�Y���'�~��\
C��{��:��
wc{0JU_��܃rH���ݠ�/#~��*� �Q�0�J�6�H�Gͤ�jA%�(�lE,-s��y�n��`�=�;���-ڒ˟J�.5��^[��������.�ˋ-5_�DxEH�SdO�w��%഼`MEw��h�V�G�D�ƙ8�fT�J�!�
 � �����8j2��Ь]�!�;Ǹ:�=�.ܘ��Ӧ:U�����j5���4�ѩR��DVm ¤���o<2N�i��U�?g�m�ݫ�zw�-���Ӳƽ��D��p�vХ��K}��<w$sh)i'�w��r/VO`�'Μ�I��V��b8��_���`�'��M��3-��l�-YY��8�'mK���;AO�c�+v$�O��6b�W+h���5���^������~��dS��W4����5��[��Qn}[p����߅��h�./M �P�*�	���3�w�HB.�mo{Go�~�����j�K���E9�BMP1��*��.��k�	�V,��p��YOjfa�����θ�|w�ݟ�@Zn�`t������+����j�N��R���/���yU��z�5;~@����B���Z�yO�=��G= � �d8w	�ɒ�z����"aT���<�l��lhoΗL�����3�@���ͻ
n|HË`���h|1�CDJepuCM�`Q�J���֕�T&��@$�r�B{,|_uB���(�=~�;er�qV��f.��{z�G�vu��;�oiN�r@$|3���K��]FR[����m�ʹC��&ٜ�.xm[.�����"��z�]�^c-�:^v��{E��0��t|V�N�58rŃ̏c!2S�;�Qb�m8�/��1��������U"�l�f�%+����U{p�1p�r����6�}��J(��]���*�@;zV8}�E�TX0��&�V��5�nt��t�O&�#��� 7�����{��ɍ&"���!7%��&Qg.�v�FhRU�4��o�q,@D�
�ޔ^G�sֱC	�!7�O�K�����<��r���9���+����e��Qg���y۽Y�U���c� ���d~ٱ�P`���{�R�f�Tz�D|��q����S[3�܋�S�\�֋�V��~f�CI���~������`8�W8���SM�?a��C�<�u�mn!Ca j� y���&����ؖ9I�`�U|�c��h�*(��5x,jH����/U��U($A�O����إ�[���% s�A��ISv2��M���?�aA�f����4��,��9)[�<��[zm��r�Ejq������E[����B��nWи��f`b�v\x���� f�x���ۛ�kMjZ�Ӎ�8�vO��K��7��̱<<�&+��;�;�g6(��f���X������Z�c܋W����u
�:�ôj:v�C�~�*!� ����>�zq������~����X�+�Ϋ�2����ls,��Hd��E �������	��S���U����Kj�P3�
�N�R~������蕅z
�+gAաfG�d!hi���Yբ��ku�{AWV��@h�Ҹ
����Zu� �����EX�M'�P��{xԗ\ji�n��&_I��O����R�t1�&l��ۤ�lD`�5�8�ёu�DH�.Pʎ=v��r�/�_����
	ْ�����j�b\��h�Z�3z�ս���?�s|d�R�eg/�T��:R�S$��N�{�˝6c8��ߓ�)8�"C��Q����*�	l}��������<�0m�P�ܑy��2���5�4�=F}EH���_(�zc��2�H� p�6+e�l��X��@gJcQ��Y��a�2�a1@��M��#���Z��Y�{����#`�UD���	f�-�4:[V`�`�kuE�+>a��k2��w!f��S���R���t��ݼ��3�
�>���B����F�Z��m�Β�C��З�s���q�/dv}�Y$��y�}'�̀Ӿ�e5�{`��C5�6�?���߽ex���o�
!�4�闍�`�,r��64Xކ�Cn���ɘ�,�G�x��
����n$�}�٥B�L�^m�����~y��D���*�=*�HҝI	^ܪ���Q�}��[E�m���߬�1�-��x�IP m��i���h#�F��C� �E����i�,~�j��)�~rE�1	P��г�;�0�]a���iQC�0
��B;}�@>�q����̊��0��`�e:4ֻG�Ե Ks_�;��m���z�`"-��s񢫅`a�g2�^�j:u���";w��҈��jx�1��ٵ$��7Uj���t��=������Vа
���[�
����y�M����i�؞6B�%���e��m�cxg~=>������;w#M��lZ��p�Z
���s�g8@�Y����RW��G�l�կI�s����f`���kz�ߒ8g6Q�6R����t����Ӌ{�.�AK �^�8�Q�� W��F�}kQ�l�	�� G��5H2~�ż�dud���Y�KhQo�l�$�nz��tO�u}؞Eq��q^�{��p�h $�Б��"�a���K�c0�ќ_S��S��,���6�#���MY����T��F��"�D���Z�a2|���Pw�-xS���c��7�&��	��P�)��p	��bO �`N��&�-�	�6�qNf�?gpN1Q��n�6+�X�Y���]4��ho�9Q�=������gX�O'�Ц��,lx4�����Ԕ덉�8ߜ ����㨫�aK}~a��	�6��l|P/��4��'���6���;�yjIA��a+�tʤjhc?�S9� x	q٫����;��Q3�g_��-[3�<�lґRZo��tx�����*	���5��גI`��Y��T'U�EAQh�M�&|6,�Z�t��`��TS�V�գA�Y<�>�Y�	!���q���E�I{�Z��.��G��i��)/�X&�x�Y墌�E��]C�	-6
�O�;�s��E!�@>�f)�>�i�M@��:��K�n���Ώ���ݿ?:+C�Ѡ���̉;���K ��ZScF���̊15[6A
�<Aa
?�f#."��(��QZ����s
�;���Q`69���j���7&�j�՗�G�Z#��j�A5@ @&��aD��*) ��湆Ϋ��?�z�~�Q]�ʹķ�4/b�d+��u�ʛw�������q�m��
�F��Q�]��m�gj{��8,���	_�Z�A��x������2�x�iY����R ����!]$-��v�_x�Q�2��0F���i�����S�C�v�8�A��I�(��n��\�إ�G��ǖ�y�kQ�Q*m�{�]dE�H�����͹��5N�Y����bՈ���~�a��Y�Q����O{�k�k��T�y\�����XG)��ڤ����5eY�𻩙��nޭd���%��~�=�_��n~�B4�A����i���H���9.�s`�AY]Y�8�cG�%�����hr�`V��4�g���������c�-�(?8)vUF�7�^�*�V�jW���ڧ�Ѫ��b�!G����Qm!�$�Z�f(֝ �G��w �+����k������F�N^ڶԥ�~�F��r���&dB����_�X~�9�
��0.�w����+[I�fv�늶8y�z%�0+���Å�	6+�q��� 5��Eκ���o3�g8J���PD��湜�<J�x�"�<���X⚪r�\�v�)�`�^:{q_���J��-�骒�V$���B�V���ߢD�]D��g?u?���Wv�İ��f@Q��6s��8�,�wi; H�h��Ie��emėȈY�g�8�b�&�j��J�h9��u#����C8��;��	�����,}rzĚ�O�ۍ�������� �����ۡ_��'n�����"Bg�����i�6��׻�\�w6ίGX��먦��%Us�mZ�қ�����E<q�W�K�aܫ�?��=9x�͚ZdRpb��n�z��9�d�s�yV2�OQ=QC�u@�9�'�軑;�&���|�D��/�v���pu4Z�?u�rлcKХ=��b����D��5�.�H����Ѡ9߮�����*(�~Ȋ3��k|�B�#�f�.~�j!�Λ�N?�"��R�@�-�@{�NB�i&#�����cW�IX"r��G4�-�=���F5���}~�40�x�{LZ˘2�PC4�̕�G���V\�˫�AE׸An�\'�6-���S708�n���W*�]Ĭ�^;�/��	�,���L:��p�C���aꥌ��X���OS6�f��a���1��/N�R.��Fy�-��{��I6s�"L����&��@���B+�ŋ��J�[�恁�~JE��'�X��Pʭ�ʬ���ț*bz�S��;J���;"F'���X�
N0MH��h���,(��v��oܫ��R+���>�"�H�9i�t�؀��e����!�n�K��`muA)����-�Ä���d�S�$�[ݒ���Y�/8ư`�+�g��A.���O�����K���8����v�jg���.%))10������#�]Q��1�}��0�,��Wv�ĭ��T^"'�_��9�*�&�Y������(����Qm�|?�Hɽ�����h��K��QA_Q9����{1޴���G�s��D�+��;��%u��r+�Uc!8�������}��ڝ58f�`��G�k��(v���R����:��q�#��$8� ���G������K�е�A	oM*V�Maa�������*A�j�[�pR��P^��^<�1je؛_}�����L\w�?���;Џ�__��e�O���P����إk{P�=�C�j&ݑ��'���P#Z�h�#�?����$�u��X̝�B�xJI��b�Q��Uy�B賜C��2��j�v��!zŲA}����~�	T^�8s�W�n���~�馬6��(^��8D}q����iwD�N!���V�S.�4)�n���]�)?�����v��?j����,R��v�J�,k
j�����y?�V,��`^<�s}�栁������ǞI�t$+�ud�{yO0>�e4����>s��;��'&)ސîAW�r�.`GD���&$.X`�r�i��_��ip�����Q��ƞ~wC��F��t�_H�o�B�R�T������J�=�1���%�=�hE |f��^�p�%w�-�
ˢgFt�Mʔ��'$��S2t|�1ߐ+7jY�K��|���w�d��T�Td�-�^����9�Vڴ��'ӗ��g���b�=���_�8	��"a� ����$G�=e�3��&��.��N�s	� -�l�?<����[V!�_?d�̰O+Y9�*c�h��)ή�W$Ԝ(S�ds
e%�Z2r����I���`{"�);�oE֭�3� X�#�uV��*��b)j�#���W����l1:2O��{�R�jK*?;z�I�1?ƙ2�k˄=��a�op@�kAB(*U/�h�|%��H1�3j��,�lJH��Ūޮ�����������~���քZ���!W�Nm.�S!q����CV���
��	�O���yz0Hd�8w�k)��=����%�*��}^��[>#N�3ȭ�"J�lZ�E�4��'���J�Έk�!E��1�F�ܵܟ���w0�_��xc܎���-f�����i��	�y2��ޅlA��'dϮ�R�P�s�j�,z���WЖ��a�un�/[3o)n�Њy_�k�p1�؃�	�:]M�+q�����+�"�B�x^H�*�:@��*d��H���=H՟�$J��$[H��ih�U�a��+ΐ-DG*U���3���f��edyPs�o# �*�UP��P@]����"�����M�4I?� � �GW��}z,�MU�+�\��:e�A��⩏�o�� _`_O'h`���~���M��5N��핬Qm��G�@ 2�f���i�l��� -{X�Z���\ie��4A���~`�ɀ�#㽝�ǃ3��1�����u�+���) ��!���9�-�DB�
I��{s���?s~�f1�n�����P�N�W� 9B��A�!`x��3QK/�.Z�$���YaS}�^KF�h߯qfa�x��%@@�[��¾V�ҙę�b	|V����>�2/[x� Ȧ���Pcy��H!�j,�Nt�e�)G�c������j�	�_}fB1�3�y�񚆔;	:�1B"��ñj�=�����Z�m�`��$?�'�\��U� �*
��%
> )�\\�E��� ��76�DNkwT��;��p^,��_dnY `I�R��!򵘿q�dЗ%��L/1�xQ��d���|�/4�ZU��0믖���ٲ��s�Vȑ�x��QG��ѹ�Т��rMO�X�\����tY���jcJ^�{K�)r�&Cd�g�N���4߬�$��xʊS	�i���!B�F�r!����`�^O<��}Y�35#�D�L�(s�C�ڣ���9W�6�$�T�Fk_��Ќ��ezU�]+|Rg|��9�<��u���%
�NǦ�g_���@�������[Q��n�sj?��q��}��.a&�JC���f�_�e���-_�,�
����j�'6��ڈũ��X���������H�K�1�7k֭��[k{OP�����mz:��F}��M�D�)��=�f�H�
�>��:��?	qf�G?nw\��M�L`��w?���2��mN��C����2��Λ(�f:(�k[�����c��:D�⚌�.�o?�������6�
z;�X����g��&ZJH37$\����!����7����]#ە���F�Zo��j����g�����/�̬ܚO�4z�����L%�k�S˱?���?2�4���r��0W��g{����yK �3>^ۗҺ>�H��-x��3�w�,v!��]��uM�Nw$ԯ.��,:etK�2���)�j���rhT�5���|�%p�`��!C��[��v����^�L�|v:n�1mb� a�z�;~S��l>LEԮn�Ӳ6=�K���SJ�w.��8L�J,�X~b���b�B���.'������0u���9_�S���6*�U���ڲSA��O������W.�#��ƪL{�Y �p�Oda����W�ܭ���\-�(���/��
���J�d��\�s��@83%�"����:\Q���#�c�qf�ՙ�v�P&Ą�
սW"�.��k�`�+�8�9bq\9�B"����?`T�#g����/��Ro����I\z�h�CJq�ZgH@�`ӆf�M	���H��Q�J1z��,����-����|���h%YU��p*eܬf�֏k�^h�KL� �kd����L���@ܞ 	
xw)ڛn�K�iC�$�ج7Z��PU���c����S�p��WPt5�����~
U+�;�F��WO���P��o�h�zG�,�Z�<)d�)>�%�m<��ViI�i�\~�T�&(
5j�X��ꄡ8���ʷ�5n!�`�Ϧ/���*z�0DH�Wb�)�;�.:��^Z��dV�',.�!��� ��>&��b�W�VU+L3����<���s�֢cӒY$��Ls&P���[u�����W<�ڇHs�k:ƹ���A�|�+ׁc�b`R%1pdhxB�f?��]װ��3�'<�kEf,a%C��|�c7��\T4�A�1l�ؽ�;nj�:�r��|�/�Ο�h<�G4;H��\8J�T�_w"x4�����g��0Λ���v&�R6E
V/0	v,��<X��L0�g�Q���}#�u 2w��ť��H�8m�q��]�F��_j��N��.�?���
#�*�s��xc��,)!5�H��U��_��I���m�~�e6=�ɓ��=Du�Ho0�>�ȓ$%��˸���b�'�>Tq�V��_������F ����A���G0ɜ�vs�Bz]@s�"mK�h@�sMo��?���L�b3���"�ξy%��n(�Hvê0���*�#��|�%��?���Oi54o�E���l����qW9�9��)�|���u_ā���X�&��؄	5����(��A-9�q�`�TaRH�F�]��ӝ?� ��`/m�����sfrW�D��F��==*��6l,A�Hs�v��Ez)�G�n����N\^,h����~�Ղ]��C'>9�!IC�/���5m��7*NW�y��ׅ9]���#+0����`Fe��ҙV/H<�{�
/�ւ�K�i=���Y/&�����
©{G+���;sw��z��к$�
�����΢���2�/���"���N�L",���_"Ǽo��j{+o�����[L��k��,@��L�-	�B�����5J��D�)�����-T�tyQO8�\%�d5?Hh2E�:Q���|k�|F�[�ԃ����l~Q쾪#=�*����}�
p����c���;͐WJ��v�)�q�#K�ȅܙ�=^�c:c\�nU��fN�"j��y�@W���ps��{R$X��8:H�H-Q�C��� ��TQa{Z���7��k1��eʙO���=��i��S�d�M/��	9��/+����X�!���fDl�#�ٔ:+bw�S��yGSĪo�����w�2���Ѐ�#EJɾaBi:��3f���������=������3�e�Q���oc�<�!�v���I�F��d�!�(4�ώ�u��"�ゕXS<;���>�)�U�j��"�c}b����?Gt�`��g����J��x}�f��[���Lu:��ʫ�`s���e�)a;^���h�Һ�Bl}���h0<1E�fW�~�̀�"[��q�q��TS�v�<�5ܙ�/� AY�⧻�^��7G��j�=j:$2p�$�;VNO��'Ϭ�!��j<^l"8�/�,}h�"DaJJT�k9ip�~�~PX/�&�CxuV�t0���#/$��J�Jʁ�j�̟ւ��*�����Ë)�ӿ�7B
�G�Z�H
N�@'�^�B�OM_o�]����"���ج���Xy��j_jԗP����8��`7�:���@�I���}ArE7 ݎN�Xš'�;RX�cK���+.��Km�����@R,�?� �&��A�$�~o�R �f�/9�0c}���r�'W"���l8����PB��N_��r�l��V�ݟ�Z���l��X��ۿfj�p�
l����߾�sDٳ����{Ÿ~����\hCV�L�Ȍ����՟��>H�h�6��Q7Mˌj9���*�м�㮺�M��L�s���KǴay�	#A�]S��SŖp5���*�9郏�wŲ|�-�(Sd���ʆ��6X֚'�����
��ѝ�Ug#+m�h�]3�A�����M�>B+��ܔRvh�����]}���W/o��dj��-Kt�p������j����є$A=C�v'�����i�&�=�a���Dt>���� �P���;�_���\���,AT�O*��S�6"2\"b���g�R�`_����Ie2K���Fse<��\0���G�}� 4��	��J�9bR/����#\��RI��ݠ�.�su&g��#��vyF�^���H����4�Ʊ[�{5�����!㏙�Cő��K���Rj���y[��ͧ�*7j���@�js������a��OQ�����%��(]`0M�f�x���� �Iۮ�׹�YX����#��#�|1/C��f���<7P�K_���s\��P����8���U�Ϫ�Җpz	���P`���q䭶i2�tZܫ�bX!p����5��$v�Ȫ'���焽���{xz�\�����uyi������Yux�������QW�{N���V�=�S��~����\�a�}�\���B��ۂ�Y �Ŭ�T&�`�8����J�?���p6mH}ϥ~�I�y����h!��P��!�x�l�φ�v_�lݰ�!�T�o�P����Č4{:�qZi�h�e�H�Rh٫��,��3�ڭgi�@7�?��P��n�35h]�� �'A���ͭUS��i�lN�.pG��Nh� LGv���t1�g��zyR� ��u����X�%U1�yJ�&&zHsީ9o����E��?\�A��?=w�+�Q�`���@����qO�����1Y��������#;��AF{gZ@B�RЈ~!�i��w�ڀ� ]ٿvLկ�h����\H�!��~����K���T���`���3��kĄXF��a.�� �%�� ]:bv��>BA�\��4��X��ε�� ��Ǳ`1zz�iG}U:L�l]2g5AЬԅ�Ly,�N�XM����n�p��d|�G?Z�l����'��y�
4�ˆ��a�@7���?�Ω�4O�P����^8huzh֛�BS�Rg��X{K�X�4	^�YW^$�q5�[��c�����E���j�[������㱼��rD0��9I��P`qzM��*�iYg1�삽�E1:,[w�-��4f�g1� T�EVU��� +jdsP�omP��X��'l�}��
hn)g��b��}��(�*�r~�4��3��K�	��DY�4+�ϖ��ݰ3!�n�gӗl/
b� �y_��"��e	!\2>��|f��uЕ��0�[w�
��'5�����Lf���1�9��RnM�z�Wd���w|�8�� SK�U�lh� ��&���岙���B��W�%J컥�_�"SAJ����i4/�t���Y|�H9��z%8�'��P�X<mu���/ �{�=���Z�e֟�8�ȞH�Ϛc�3���4�b�q\E[�ƯTŗ;8��Cc�<h�������W�a�
�Ӷ�NpD[������Ld�P���)jd�#�E��}>��&�-1��Y��˅������̔|�~@����}΃hң��0�S��n�	��W�&W�	'���Fe���8��c�7n4��P%LT�O�9\nf�~�}˵t���r4a��w1xh��5���pe��pYʆ4��	d�k��l�1H�YE"�y<���~;N�p᳐�gW�����b�vGU����H@_0��_N�`[�"B��z3����hZ���B��h[uӒw�Oy�ߜ� \�E	^V��_�����Y����/�TŇb�G�+�Zy̧bOY��C99�E����P���v6��)�ڝD.|��j�ǖIY]yG����gu�������?��s`aX�90g�tE��3V6�A$�n#c+���9�˭���[��!T����p���-���V.�!4W;R�C3�[�<�-�w���v�0�S5H�i!�HMb�@]\�x�x �2J�Jy�!;B̾�L��MHU��
Q�k e�)}/�W�'W��o���%O�,��S��Dz���SxR^a�)�8�v1�B$�}����������\��&y܃���I�<�?�_Ji�򥑥��������҃tÇ/�
����-Z���ΛhN�|R��
��"�����3����ËCz1W�#x, K��.l��o��T� 8E�� �Wd4����[o��|��A��#E.�-y�??��J�Ү���Nyz?�^�|���������<���/B�(�}(C�.�v�e�5���!p��h=J^��*�B�P:<�j��M�R�̈�|C۔g@�X;f�f0�B{��%}W'?���|�[����k!y6��l@�4)ы^�����d�R��\�8N���#���{�NǱvV�Z��`^���Z��f��?e/�J�J`8��iE[�s�.'����Eô�C�:y�E��*��T7�%i�-S�,���.���S�B�gn$�:8*.tG1��[,�H6�H�m��~�ӎ��D�^]Up�S�)]�MFGv!�.������w�G���T�i5{���J ��D��J+:Nfg��Q���dK�~�.�>*�r����1��S�#tU,��Np�ѕqb�fR��^N��Q@J�z���ϱ�|-|�[�V�@O�eC��r�͹t�A��Dr��9�Y��t��4��uiyP!7�n���pH����I�l�AG��^.�)��$�I�B�^���P�U��*M;$� 7�D_bg���(�J� �]�4�k��|�m�Aj���Hl���W�G%��u#��[,G��4{"������? bN���9�9��Lr�Ì��v���/u���2�/�"��7%�%3 ����%@�i2���H �r�~�Ngft�z)�60E�n���H��L�Ŝ��]����f^�C R}������˪��Hl�Ob�X���S�=�"�[q�?���z�����/�Zt���Q_���N�K�>�{���"�3��3������������?�ۼ�_-U�C�B��ؖ�����bf���?���Uu��k��KsL��1��0�"@�DDp�	�9��	�'�:&.��t��:�~bj�e���xCD�ʲ�omO�n?�!V��J�2�}���� 	��"�f��~��� 6�#��s9�)�i�&����\�'�GK5%+�uF��>&f�^�.Wh�,3|��mԞqD�JZŧ�ד�x#��x:���h�Dh{>�ФS��+7���'�0<�(�J֖�QMR�(����Z�c�"?���L�Wq��Ť­�wfs�V���Ȯ	
����W�d�N�L$pt5�n����6��DNA�����N::~�{�4s�?mÍ�M%㫿,�I����bjD6�(ˍ�V�
�+��H▘#�7 �qz�Q7�v^LZZq��|5
*}y��7��9�c���7r}�b�����2 ���P��$%xk9������>���%�&����@Ą��I�gq"R�����gP�ܔ���H��S����	5<b�m���3Sӕ��wa��Ĩ�1왣����.Q��.r�z��3��bSJ�<�1;���5;"n/?���=cA�3[�5	�u�m�2N����r XMt�$dJ;}��fJS��9�{#,�r��ksy�ߦ��@}�[W���D�L�9�
"�ݼh�HR����x�? >���,�Q0t&F�E@��5��`k��k���rPm���ni��â�Li��<�����rL�ob��xx��k(���;^�F�/�|z�̥N[G�Ԣ��;�Z�sG7���2�x�l�,#�D�1�[Y��Hi&��)�xJ���F0*I����w��?�!۷+5�N&��d.�
�{�h�G�7���魺�P#�Ұh���rŀߜOϡBQQ:-?zm%+w���e�����ՐĖ�;�+�sa�%�[
�g�Gi
yI�<)����=�1&}ae���Xd����t(�tXA=Pbۑf�L<*��p�_Ԋ���P�3���$_ts.�#u��R�d��7B���XH=[3B���� P2�}��,�?����p3��_P|O �
�1�d�S~�B.�u�����NP'<��K�K�rQ��@�V�S�7)h���?\��uz_��[�9H�G7ź�݈"�05������$o @7xu�nPm�5DB�~�Պ����7���}���1�G�R04�e�Cb��%�t�S�]&��a�1�4zݴ5���Ί��.�7%���u=*��t�jp!PԆ��qG5�I�lQ�O�����9�lY)��ӱ#�ilVu������3@q�
�}8ڋ��m�&�(���9�0��ZPI�������0���^2͔�֮TkѣDb�_�r��"Ee��<aJ����Y��'�2U]����䷮�q0�u/T!CA�'g�;�Ȯ|B�u8U[�>�rW�lE����U����_���S��Fs��`���l0Y�S�M܍�6�Rʬ�ʧ�7܁g����=���x͎���[��VL%f�t����7VŨ�	ąQ��^�6AX5_��#�X�|5)��k��`Ŧ���1�sA<���V���2֤ܫѵ>)qȝҸ�k�&�6k^dħ��7I�&qv#��%�@_�6�3W�@��&�~ډsz�B��")T2TE���s�tAõ��� �{�O��� 9��I�#>��u�bdp��{E��F����e�<��4p�^ŌFBQqRe�N n(�f|�F�%����;%W�~�AVb�%�9��1g�0�?(�LL`��U&����'=8uV_.�P�STad��\h�R��߉Mu�taC,8�}�)�:�y.�@T�}]�]0Ջ)3Z�1K��t��I�TR6����ڌ͇α��p	Uf���>���Uʆ`�m�֟�3����#j�����'HJ�'
S�ɞ'M�������د��n�ɏ����TE����h��|�K_�-�yBRc!���G�+��+�x��'"��2�m��M��)�S�K�����JJX�h�o�F}�XF� Ȫ����q%�q�n^� �f�ʐ0�mFFj�F[v_���w��=Hd����t���1�{ �]X�0�Q1?^D�A�=L�9�����g�Qq��{i���G_�ڌẓ�ʆ�M�O��-w?��t�y;yђ\�f,Jy΃�*� B��R��B/I���-_̌i;x8<,�%�)��ӻ��F�$|)̌�Dh�m�"��]�@�����r��ǛS���[��I��A��8�i�JSՔ��Q-_��u-��%���'����ބ8^��;�����3���{n�����ռ~*��X@��v������;�~=u/j,�I�D����H���8m&o�-BL��n5;/`(���VB���lZ<����kG%�D&�$
�W��?�nxX����J���`��Z�EĬ޵R�E�۔�A������v�y��>��R3����k���BK`2ӑ�N��i�菹�y.gm�ˊ`p8	f�������Ғ[��J��lW0Bh�����t�ͱ�&���(<3Iu8?7aP�*��햞t �6Ӧ�������GZ2:}Gs�.��i�DQ�i����)�r~���/8KK���A�DI���:��k��� �?ahZ��P�����R�l&z`tmj�KE_�]ƞw�]F����q��??^�UH U#�v�W�� �=�ΐ,t�7qlh�G�W	��)�w]�|f�ѹ�3�'s�֎aa��C"�`��n삳k�-\�d(���H�Րho�+���yͪjR������y�"�R��3�R���׃!���gs�&q�k�
�:�X�0�?9�4=x?D=� f0�x<a|��z����O�4Ro[�:o[*����xvnĺ)N��٨��g�PL��vbS+!t���6��,�݅��2��+T�J����k5.�<��qpx7��ީ������)%���09�,FauJ�[��P��'l�Cc��N2�s̞F����ǐ���Z����+de�O�����ܽ� �s-��0��Z:�B��Ёk�+�N��Ҭ/�"���b�� fN2RZc'<��H���^7�wQ�����F��lṘ� w8����']�m���Ai���� 1<X89�{��w�/� R�ށp19H{~����ڎ�WW�mJ�j"ZmQ�}p��'
}c�c6@��$��K�9�e�@P���ௌ+AEo���A�ݷ}>$^"���� o,-\Fy�n�uH�\���QeS!S5����0�9�IF~�xg�?�p�g۹i�2+�
kH� K��'�!SF��d>�̈�ؑ��Ct,�P���33���˴�s�˝x�Ӱڏ�pt�7�h���ܯzp?[q����d��
ܝ���d��ZEGI�M�v��-�y������Їӄ�Gh�L����̏Z}�R��8��QQ�=$��qv�,b������T8��T��("7"�t�ףP�S�8O�T����<1
�����/�Oq=���Y��T�ȶ �H
xnX	��S� ��ͭ����R�雸�s�z7<���R8��D+���-�1��l�5�Q������HsFvZ�A6@���2��B���V��za�6���#�9�(���OM7���W:�x�k�߆;_���I3�y��e��@��'���K ���:�ʋ�c�WLؓ��w9�������u OM�)���.ŋd|(�E�~�$�L!qP	j��M,F�}THJ4���I�U;��to;HFĘ_-a0�T0)�Ь��"�	6l�ExI��Ң_�6=ip��>�)6��+,̾��	[u�a.}]o|����Z�}��<9)�����H�=�x$R�Ζ3�U��19
d�o%���<J�V��t�#�WҔ�.]��L�bv:'��O�Nm�`�"���F4H��r�3�1eJ�T�z�|y�'G�z��U`M��"������BE�4����Y�:i�s�H>l_�ľ�2��YT�6?;�^u�]�}%��>�F���H�G|<F�J�$�~�����%�I� -���L+�K4���Ҩ� G��}i����	O��;�rG�(���v@9��
�.
�9�E-j{$�L��憋��"Zy��@��K�e�R{��L���Z�9ǂ���
��$���O-�4�Jv�{����@�8^lƱ��M�!�6��O&S�I�@�������Ay�.;kXz�{{�)���vr�Ah0z�gH����5N��f]�a���j�n@w�{�w��4W�FR��Ks�Wa<�mlS���6<�����ə'=��n���'�6���%���B� ���gP��Cq3����FS����X�?;�vC`~��#�=��rC<1��y����O����~����0��bܸ�l��L�P�F�Z� x��Z+5"�BaNDy�"�]5E^y��)f"GZz�s3(����Z�Ev���1��9-��x���T�v���,4�Gíz�d�՗/Y���0�ʛ"ˀ���'�_�ݳc&)U:����f^��Q�u����0���
(�dD��͋ޮM�rQ��T(���}R��J��ݺM�5��c��]��G��6>ݯ^����@LMg�y̖����y��v��xWhr�ԃ����5��V��<����vxdռ��zn��#��33<X/i�b�K� 
�íz�RM�K����b�n�0b=���mi�f3�´r���g
��Vx�v�[���g9�i���U�	C��XW�u���|?���D���J�ܰ9��&y���A�(ie"4�7G�c�Fђ*&���K�to�&6�X/
@~oχwMa��w��t$�`�ߢe*������+(�$o{p�T ��;�i�p���

��|�ޥ�����z�O��w2�Q���9�i`�
u�n�P���O�Va�~x�|������8SVu�J<P�-���%�\gԆ.� �_������^
HR����rĵ_'E������ }\,`S�'�v}튵|ib&p�mq��1׀����3�0`wJq�yx&�sr<(�Ϡ*B��&���:����T�[|(�K.I3����CV�+@����ru>!�|�"!�\�l���KW UMy��j���?��R߄O��M}*̤�~�jrϼ�(d���)���<LE�T,��I;�sn��.�VP�d�=_���J �䶨��܂R�b.ͱ�Mh�c��&SJ���ft�u�z�COL"� ��Gx��m`t9Q�k�_N���T�v�o/�U/L������vd�����ro���v<#qU	�jh%=\�\�����}�Gh�^�5H�g��P��$���}z�UP�� �uc�@2���ê����̜mI�@�P���= �T<��cz������W�����/gbp������n���$X��η���I��8p����x .s�-�:�@&PphC��tR4��2�"���baBr\���(��O�nR�����20�DV�|�{�.������}�Q�u1���=�V2/�h�]gs����p)h�L��B
�inn��r1P^.�z�(k�H��3�Ub�ADl�?���~D^����{>[������3�a��rC#/�J����U��#�������/9d,����+[%����v�ҘW5�gz��׵�d�
Ϫ�2���`�_�E*]�����T)*�Q²4(r�1�L��~�C>��6��kp�1pE����&S��϶<�]�
VY�gN	IeI�K�"=��m�(ѕQ
�.�%�P�M�p�U��b_C/��Bϼ�I�L��\0��⫖K�[T�
�ڋ���N�֔������Ѕ�t�J[T	����oԒ���d�R�c�˄�]e�a�}����0A�} {�T�౳�nމ�E��1SC�ᬓ����\�Ӯ\�a/�4'�]5��	�0���aMj}��A~�賻�y%'0�1Zs�@cK�Rn��L\>��KP]a�>��X~���9�����'��{����cɠU�|Y�CA>��Îg�������У��_����e���eWd�5`o��+ʭĩ��1-�q��?�$��LNQ�>Z��ģf��zg�O�d���n)��?Ϡ�f`�����#,�BI9rB��J:m��D�� d��m}հώ F��W7��^���W\��;���[��,ޖ�r2Q��;����S��)�Q]%�9js�?�0����,Ĩ41|��X�I�tP�Y&+��	��K\s���M�g#�����'5�,N�J�R��e��/:���*5H4
�W�^�2PO��K(j�	��(���zo�����6w�'�3��'�\ј��5�/<¢^
�O��/�QG�"z��I�����lP57�U�z�"4���[�_i%�{�}O����Y�l{ ��Y��?Xk�a�iތ��@��q@D���isÔ�^nڂ�a�o�h����k�j�Lj4�3�׾5�N�Ό��B>Vx��W�I��d�]����쯅1��
�6�}Y�{���
����#%��Ca�
����7rI��Y9��`�x7�3߯p�� J�?#c�#��ܦ8��!�C�(`0�G�8�#}���y��Y�\
���q�����{�ÀW�A�M�v0ұ�;���A�Î����ح]r� n�G��g%նT�[9yK���J��xrFѨ�k|��S��C�*N.�rD�����	+��%�_�H�G*挰�>����QS����+<���j�O�/
~�`��l�D�<}8Q�h'��cp�t�c�W5gV�RD�BʫȦ�?��2��"ڜlF�ă)������=�-�	�ϸ��0�Y��*J���\��ԏ�V3^z���f��#ً7( ����юh��`�a�jQ���u�;����,tK5;���|�2�I�@����)nr=�Dv% k_�%�$�Jm�s!>��{M��:Ԕ��W��ֶJ�h\�(�(��U�@�U1.�T��9.�����
jY����C�B
*f��� 5��@x��L�r��+O����I�#�z+�Ud�r��"[0]6�Ur�^�'�|��@���]KQ����&`��X����A\���J��������>��S��N}�Xk�9eJcGSW��^u��shQ^����5�?Ǘ����K�o�Ɋ��t!�^�X�,��ٟ���b��s@4J[vo����^�m�V�*�w^r6��L�� ��W�������vD�y��1�K���V�.0�AAl�2�E�R>Ȝ����G��� �/�?z%%��i�&\^f���x����ٶ�6��,Z�����7yf2
������a3{b� %�<���Q����?'�X�p�<�!�5�?'��3zJ,ɧ-bW�{�M��e�x�E�C�P�Y�@���2b{:��b^��`wBM�9*�q����܈���MB~5�wa�mm,��h�T	E�ns����Et����wst�MӨx��i�h�-z��z�3�D)�x�ahi
��j	ne�#	�S�F��&�Z���l�uP��e�m]�4,��;�t��|��"z��9��f*�~-��j&��n��"l��C��N���~�2�>�@��)�mxh?��f���B��$��ꊿ���]7�D�I�Gӗq	�*Ьڢ��i���A�A����� ��	s8�+DYY����ҷ�_��~r�c=Z������6��J�?{oVOS�*q[��x�?��R��lٰ�vϞ����!FS|ӡ74�Y����[�^�d�������7�~BnvR�خ��SPBr�1�J㟲����\��PK�i�')*$q����#�_N5Գ)?2C�����ĺ�Bl%��Q��ǿ�CZ"<L��_���P�ŉ6�� :�	iP�]|XId��[��蝾u/wȅ�٢-�[��r�-��g�T�h��e{e��^k�pLIS�ytE7��C��J�=�����_�5Mc��Z6ƶf:���� G)��7�!�q#�n�}�^�U�`�k��}��C&��ѵo9��10Z�s|�x�m�s�%�(Pb!����f��p7[p2�,j�Oֿ�^���ٽ�:<@�`�@��'�p�À��x�K�v�������u���kX�S`hիE��L=���pOI�@%-}*T�������&��a����*��q=4������J}2�I�kĴ�v:�Îx�"��Y�n�#�Gu|H?�������Nc�9�� ����Dg�K��B�^8��I��S��}�X �y4�W�$ܽ/�M\e�q�<��&�L-/��Zn�b�:��2����1'� �<��U�o�w2�����uE	�\BMZ��_d���T��:7�$����%��U�߻W����DN	;g�B�؄�0��k{AMHt7�+I�7�pu03�ް� ���@�#��k/ۇ���$Y�ļ�2�@I�NC��,P���Zn�֘����� g���s���uĺ�Q�KtON�La_�@�*
-��%7��M��h���P�)�
n��m�F��4�&`c�ȹ��wI�f��R���?E��Ɋ��s�LS�/D1�P���w��� �Z]W5>�� �D���Ux���\�kLE'x���DP���ˑ��RЖBu�!�W��C�|��X�.�g�Q�p9+ˢߑbl�����M���h���z��>	l1x;28T����[������w���z����"/EByɈ��#H��ef4���ˀeT�f�԰����=��`�,���#�����w݅	�ם��N#��b#AG:�_(6��/*r�󗓑��,6���8�B�=�Y�.A`D߄V���燕ط-7)�j���,�� ���3�n��~��,n͏�=^ڟmЄ�� �B��"��S���!qۓ�Pا1;�j�>�)~��x�0:������"j�)��6(�S����w����L�z+��O�n�a�:�=̠xw���+xw|eBr��ndi�@��b���N)��Mi���wG6��gK?m)!v�.`m�v�r7���ժ�6V?2,Pk���jNr��ϛ��p��44rQ�KlQ�i򱳊R���&`�����l���z:�P@莒#���ғ
l �zo��Ӱ���ǇU���IT7�ii��$�1���-�J&d�ѧA3W�䬗�_���ơ�*��C��X���q%���<�*?3e9�|�����.8�86�u���S��-��5B��!�c-:qS�5+�D6O^�Cr��F�v���,�1��}޸��b��܏� ��M���g�ʷ�YV�j�����A	;�FV�qՍ'�X���9�\�$�?�C�P+�l��m�L&e���o�;H��AB�dz3)r�Zzkċ��i���P|�|cUr�auH�kr�:���)�Jer�Im�
+��N�R�¨�Ok�Nb�c�Br�mG��>ʁ��!����B��B�d��}��ҳ��Nl����y�9S��g�|���XHl���9�n�����t��i���}�fK��3h�5�؆ɱ�J���Υ���A��-��_�X��X�O�q2��U�<�[�>`�^X�왲���.N��Q}胦�4,EL���6��UX��U�����o��Qܞ/a�2��lDg)�ܛM�"�t�:�p�S��sQ�3��BI�y?/~M\�Y�!�+�.}��b���X��"�D~x3���ug{�v�(������^�2�9C�>���P�Y:&���}����Y{� g@OK[��*g�d:��?�S��m���#&�[�K>!ڒ��{O�Nu�nJ�"�T�N}��5rE��'tE_��Fsђ#F����l�,Ɨ�� b��nB�*���mVYLu�~�Hh����^�Zh��Qs#���˦'_�pJ��us�"�i )�J�!���WiN\�2Єh
o�{�����N^H�+��l��8eN=���j}g/��gv+�� Si85��;��nK���A�I��[TbsY�)<��D�,�������>��:rF� ��o*\��x��ۓ��6c��T8�. �\�)W�$%xygGz0�i��妸Y��b�
Cp�U�95�BUsq�����8��;���(�C���6LoĤk�+���17���8�p!��rJ5�S���l_�ԝ���^��Q�p��\n�T� �z#F9�)s?[�X�Hʣ,�R�V̫���Kڥs�xRow#I��� gp�Y4:����c��k������r��S׷~%@���4��y�F��q���Vpˁ#u���f�
����:�F=e�(N���z챿���+^�B�y��%�ld���U]�l�Ē�x�iq�/1��ChZ+u�+��i��B���Ei�%�5=�,�7݈ڥT4u�+��'��O ަ�/o"+YPʰ��|yYj��>WZ�:Ekզ�+K�n=F�E�
�����&'��HQT-rK>��{$[p�$�ŭ�qȟ��]U;����r
�y�D�������bz�1������t�YFA��O%�n$±���I�+ e�`������ɤ9ܿ�4Z@:v{8�%�t�rQyK���>uCO��U`�?пR�cjB[J�!JGs�{�6�2C�!�X�7à���@M�&�d��s���B����lH��)`S��ٺ�|�+�J��B"@����'7�L���^X���.�Q�[� ��g����"�%?��Տ*��oc��:��2���C�,�y.��M�}�(P��}���̶������潢�kpk/���F]��aXbq��Z�;��\%�lM��1�C�)��c6~1��4o�������i���C��\��S�?^��Υ��w9�c��S��=����K.���&���?�2��E�R��S�Nb�}[ߢ�|+9K��2�L0�g���TH�*T��b ?����Y0Hר�(����S����a%�u���5I�Zv��[�?K�mٓA���}�U��p�5R��e'f��8���TG�+7"�<h��ٻy�Ѕ3��9�����.�/
�
W}�|>�J��:yz�5��g�H�Œ���G7�[/�̟���7&1����m����X ��,L���7]	��6E��3�I��>���4-�.�JgQ)>.���#�_`@�xe?nQ�Mk�ȕ��9��V
	�=���<J��D`q��~Iyt\d,�g���ٌIN�ͽk0�7�BO)=Y�v�>9�$|zXpj��%*����͑�z��k�����t~}+ً�p��qL����k�}�J%j�����1���l�,{oP7'���*�W�������.	�A������S��9���ʽ��{؄!����N��E~CCܵAP%�]�ϛ 9�2�v����dx�)�ȟ��`���~�-$o���$Ғ9s�J9]<��y�k�%��/o�.17�������p��H,Q�C������Kk��D����Pp�?SjB��x$R	�MD87�ͷL桨o�(�	|j6�E��"�������y����qq$�eMl�*mf�vn��@�L!�picE����~��o;�v�Fωz1]�Z!�|i�>wP�/�|���5�q Z�^
_�3��|�����> �2�z�V��ݏ��|�T�od��"���!_���@|J&��>_X)�/����z.�K��a���Q�;Ug����ggP�y���{]�պ�rss���#��Av���t`+,:��X>��D��C���G,�eiV��N���]�2C\;�-,��	�Z�F�!�h��HB��.ߜY3k�
�b	NS$4T?Y���B�"w�+��n_�:��o�4�(+�u��7���5�=b#�,�oΗR�$e��q-3$��y�?��W� /��7�i�I@h��\)T��X��
��l�3���)T!2&��3�������ar8���W�@�y%��f8��&���""]o?��"I�!��<��J`*#����i���&����p�0�X(�CeG�'}N�+ s ���#�|�B!�7@`�A���D��>����.8���0b���h8�8�>!ٚ��{B�J�9<��cג/1.�"V�df�$�{U���Jх&�[/�Av��� �tW��6��$�E����+|�*���d�c|�@�^s����7�9�h�c��;w��d���FM	�š�S��r�'���J~h8*���N��<ּ�g/��~�ԁF�dB%�v��ߵ��j~��
1�t �]�����@O�Jq!B��^�j��G5����ύr;��a�m��=�YA&���)���Q[��F�!\��f��A�P��D�����6ߠ�슘3縢 $�?r�
��O��Ҹ��O�"d޸����#j����p�ܰ]���T�䯳L����e�a4�;�e�[�*������	D7e��f05p��[6gK��r��U;Nf�{ʍ@cb��5���!j0��J�����G���	�։��k6���1J:C:؏}=��V�6�"��e���g̼�1.�J)Y���i���ۻ:9�1�����?�̗^2��%ț���H�6 sl��dz���R�/�P��?&�VXT��l�M�B+������l�cO�x���;(��N���N�/�5��g�U�����d2��CФ`Z�6����ٯ��YT�@�j1����"^�i1��ۭM�44x�f�}]f}��r�x*�[�g�C{�����Y�>O���	Tc��Wj�x}5�[%
P�j"-�I�]����礭Iv��Ռ���]X�6����a(^�I�:�Nܽ�e)D%?9jY6ԟ$v$>S}��N ���e�e��}U��f~��i",~�d�������q}5�㛛)}��|�����!���.�f�o=c���|�R�}��w��o�(�R�0l���^%l��]I������n2�*~+��7(�Pz���54H�i�f���R�r8o����Ttʹ��.��w_������HP+iIߚ���2P������-q�xLĴ-m��� ���u�[C-��(���SȮ�(_N�V��S^]+���<m�FvY1ڞ�,T.~q�"]@JJ�|�����rq�]�Õ�[>�wy��lb���,f���1����q?CV|A����y�K�(^&cU����,e(�JYCV��h�hk�>�^.5�����&��G�z,t9K�5����V�(����}g�
�fn
����!yrr��Q-5���ary`��b�\v�c�Gq�觲K��n(�,�n�r�W0�'	}U�{��m�"tǭs�tpC��C�"4�k"�S���_���۽N㑈:T�S{ѝ[q�㫽V���U���j1t��p�m�2w�mTԒ�&�����WK)���#���� %��@��3���9�P����>\�Mxd��ҎtJ/��-�����[$���������4|��ޒ�W���� �)p��D!�$v��q�6jDO��<1�������`�6�\,�ӓ�ǟ؉�=�|2f���rRQ*��u^���''��~��-?�C��"4h�5��� ��JaZB�J�aAE�����>䑒E�E���?uP�O�
��3h���[Yή�d����"r�>��:���ѵ�f-�5t�Q��P~1�<���*���5��c�!$QvԌډ�3�!��P������ږ&��ǋ�4q`��H	���S 'xy'���M!o��",��,�iY�#$��F}R6<�>�E�GA 꺁�'��zoC�J�H���b<9~����=i|+(a��:�'}�O�!Fz�뭁)�#"�@?���&u��w=��&�n�4�����P��T���<V)���OOw�{�֠st,��0W�_g����B�uXFN�U�F6����/~a�"��ȭH^���e�Q�P�P��_<�+R��'�ǎ^$�/uIt��^�l�����J'�$����4v4_3 �0�gr�4�'K=���͐��Sؖ��3���@w���M����Y�������.��y���Z��&��������u	1�Ք���s�T�_6+h�"�yc�v�z�Z��8$Ɩ�}�y-�=��u?&ED1M��r�Xv���e���lHKn9��q�����m����FI����cXX���L��1?xz�aZ�k^nd�G��m���(t����$���`>|���� o��3�;l�9�Kz^�ϲ�$B}]"}K�����Ѹ�u}��z*��_�n/p`�'�#"]%2rN�v�|��dt�j���M̈́D�e��񔴣9�o��V�+�2*u���DlUEv�N������Kڝ��a�n�����_b/�#Ag�� <p�讼S[&S�C�e?]��|±�U蔩𳌭�{%��3�ʝ�K=���LnaH��$�������j�g&��������|�G�l;��MO��G��1v{��@q�
b���w��%�P�"�!�&��ͬ���X�8g���髁��ø��5�-�iҭ����k*4%R��D�e9y}6��nZA)���t�[��MroX��P&+�GJr4^-GA?��;���N)-|�q/�����;_���Ԣ���1���lb�.-���d��엳���!��ɏ�×w���˔vh3�[��2�{�C^ �����a���~!ܺ��Z������r�~�nkp�jz���v7�/���(�� �.��z�SciN�T�'8�W�Ғ�DϦۤj&R*�������n@/�/������^yg�X���Y�X����Z�R�4���>w-��i~_{����;9��Hg��`��a�6e�Yma�KQwz~T����6	��EjM����9��^����ṖH��=�����_��-��Q9��򤊦Ղ��ӄ��6���[�҅��@{�a.x(&�C���Fcz_L�2�r:(�� �>a懆�	y@����t򑉰�_���LCa��\���y��R$���T����G��Ԇ Ne
��f?Yޓ�s�4���E����t}�U���^��K3����nN8�co�Th��`*�to=����I�+� |���&��.�@���p笩�i�1�
؞�C*'�m��A�q�.b���l��
[:�7�8i���4b�T`����bx���d��?hF��#�5X��1�"ɫKIU����a������
�O��ӟ|�W*/j�V-0�=�-��d����>c5����v���Ϭ��D��ѐR���teB�p�$�1r��j������)g����_�t��(����N�a��ٚ���2�o�?���p3��i���Ve�� <|	9	.$�Bw*��b��=����Y9�L�@��q۪�֤�Ż�B��h�?�ΙL�a�$�7-�R#Dz"�.|�"��b8�&�Tog+��X؊L�H3E��}J:@G�f	� 
m銱x&�:�e �eN��u�� ����s��0�]��_=�1W.y�,���3���'k.��踠�{ w�Stf`�R?��X�2�.�'u���<1V�>?b2wW�T�Dէ��	?vMB?
+DF�ҋW�S���@Q�<>�0��8~�!��n$���e���jh
�����e�xސ��|�$Pf�<��w�t�v��J9[.�>����g6AZ!h��#�ox�l��'_�?j(8?��Hc��	S8��Zzg���%�!O?$����t�������X0e_�8������v|D�e����Cf�^&�sQ�#_{�,��������(	������KV�	�u���2�/�޹%�P�>�l8)����`Ã;��J(,191w �73�_�cg�]�pD_��dHH\/�F�i��u����2`"�;��a�կ|�2˼�F�J� ��{K�����h֣!�,��ΒS)��p�࠲�#�͋8ҍ����^̣��~�Xhr�cz���Q^SҟE��Dna<=�)�J�H��:�X=��i۴�1dݡk���"T2a�H�{�Z�$̬3Vnwr(�\ ��\E�QG�o�֩��I��c�-=,�"	�ʓ�	2����*P�V�w����R��4[��X���1�l�r�X����p�|�1ڙ��S��ի��.a꾪��km��n(i�5$�Y�rcQ���N�E�� ����Ѵ�oE��G�K���\Yp�X��4B�wJ~�o���^�T�����rT�f��ؾD��,1 V�<M*�Fc�;1���m��W8��:�)������4��-�-�0��I(���ץ���ԩ��P~w�-{�Y��W8E��t�H9R���`���3��X'�/�F���FZ�|*��	9'wCF��i��	��SDo��]H["�u}-ʳ� 6�1�����{b��������b�����ˋH�́բs��*)FlW9p̘u�!���lu}�O,+며������Pk������v�p���g�s�Ji�+j�rJ�"Np8<�X��qe>�<����y�h�8f�������q�����҄�M�6h�T_Ѽo�4=ac9<X&����Y���±�/Xh4��`S���l�KP�1i�ۂ��S� #��a���q�����\[k@Vs�����ۿ�D���9/'����z�X��ղ� 2�F��|����u���@�`r�rЎ2o刖0�ck̩�� 	J���g��Y<L�G�J J��c������|�7z���S0Y�.@JFK����Lx��G��)BǶ�����2L�Ki"�V��%X����?#����_�p`�j�Ot��ҤP�Y������:-�o���Y����5�����!��Wq�'PI4M�	%����r�#�������/���	8K"njŊD�8�I)�t�2�����,��be����>@�Ɓ��r`h��^�<t=`�&�üm��*�bHZ Kh'}a�/	��Z�����J1�����L2/�v�#l�I�iH���ӈ�?�;���*�iu�y�`�6Z:n��o�5���#$T[/��p��i 8��'U������K�+�vUi��UP}j�i�ē�#�h>�pMZ4<���ȴ�J���h$�X�O�EZ���r�5�-�Q��p��?�k��Sۂ[dV����N�����bxv��
7>'��%��*i�t�"Yg�Au�x����MĎ�9���F
�|>)�Y�"3?���t��9I���/[yR)Ĕw`q�2�t����4������a�����r�|�8��*|3� �}��_����#�<i��|� |{��S	DmCrt�nۖ�J�x�㎝jc��Â���e�9~=����`v����ٴ~�}�~�,�^P�+Y�B���u����q�)>˗R���顰#L����5P�$�:��pn��֟M�]�:��/S�,�?XFΆ09s�Žl��X�����q�Ϗȡ-���e�F���uE%]�.��Fr��5�/�hw�J�:8�7ED� �}T���$� �(�9��}��s�m���ؚ A�&@LW�/7�m�Z�c���Ƽ[�O��f짵�G����ݤ��_}����uo�����"����P�6�����&��$�	�ԹW��8T��k��YۍF'A)��YN"�ow�A�oȦ��m�	�ۂ���WH��5�Y�y��ì���/��M(Ǭa0�F_M`�6�Aq���i���cc:�q���Ƨ�ӫ��F�l*�AfCG��@��;� �0�<批�>0S뤽v�L����c'I��&m(�tp��)�qn�v��ze}ؑ|�j�l5}=,ˬ4FK���O�4�-�kT��I˓��Ҭ�j�ox2� �BDB��h-��z6��D+FP�٠\{�8�Ż���e8�#F���'T�K*�NR��T��:��2��ԫ��ǎg��{����M;ŕl�l�zÁv�-wC�l���\�uq������'v�m֘v�g�h����+��d@i��J>MeQ�j�s0`78/�c���-C('	�T:o-��5S�O.����G-�E��Dp;%��B�,�D&�Ee7K`����R��;%�����YjS��T/j�1֕p��Z�A/��廧2°Ӭ�����Ӊr�\�1��Z
���	��t��$�.��T�4qV��\R7�Dx-�Ήjuአp�5�]5~�p �b�s�
y"r黼aή��gGY,̨��nB"Ҹ��e�"|*�}7�b��ļ|Ї'$gf��Ic�Č�S�>�V�6��:���.v�.����Ր��w�?�P�iP#����V4���	e6�����cPq���3�6�Rޡ�{��M��A2�L~Mٟ�*T�{�!���k4�n`��^���o��2�lG����!іz8��ʰ�@nC6 L@���.���OJ*�Ґ1�%=*���W�6dt��/-=�pI�z."����6�M��Lm�ࡄ�-�@Y��pT��n,2vHߗ��B�)��.$�"���	�!*���T2(zK����� �.�N��d
7�<<���/���8ٌyŤ�r�T��y��f[�N,*��o�4���7�O������MW�R��՚��Xi ����bz��;~��]l����ϒwRV��dY<Қ�U�j�D��r$��,75*�X�4�Y�Щ��k���*��7�SZ2/�L��` �z�����7������Sp�i8o��R�4$˨�
zjR	�-�>�(���vj��l��"�Z�"`���Ȍb��8;
�E�
���o_X8�kJ\�H
�
�n�NI2ܞM�k�5�r����X?�}r-�P�uw.��΄�k�i����hsL�'<�v���T(Y�a�� ���%�'K�$�/4NY���ʡ�?��'T�d]�������4oP�$��m�ẌƳp�a���(�w��h�FfR��8�U��!)�!��+��$kꓨc�7?�6������9j�-mQp+�͋��'uS<IV������R��+U@�&G�%��D�p`��q8�1�Q �,�!�C:+����}��
}���S��9�J�̝���d��wÖ&ƀK3�N:��ց��y���'��K��.0o�Of}28�qvi{�D���ظ�i�uw*l�r�ƃO�����Z�XO��!X�m��I;�Z1���6�%W=�T��Ł����O���\�s����HG�8����jЀK����}���Kb�˙7,�l��:�Xk��DkC�x&t�}B"���r��/�X����lF�#�k�c��xAi��s/�jc_�>������/RN�|<c��׌)]�7?�Ѥ�E�ɣ��a�����
����_���W�����䣋+����o��f�[*d�dcx3���?�{��,�a����k+ ����9t�0�[�R����� M�5����OC �^���"'�b��\h+��S�Η%�����0� %��o9��5Z��C@I� ¯�����W�� hbȼ7l�%EˌR�6K� �v"����g7�v��g�\�n�(j����E�-��oA���+Cz��p#��3�
�3�9��b�(� ��9S�M�K���׍�;�Z�
������\[�����j�?)�bݵ��F�X��O��%6����<掰c�g�]��E&��71��V��^��7���M*�Z[GV��2���D�'��ʀ&�$�c+��\���Rn�X���A�t�ӳ{]D��X��V��1m���a�"�8:�Q��#�c���5+����r'Z�VO+��TV��P5���4��W��P`�� �,���+���u�"�=�,��a����J	���.�	]yf=W����r�*?�ujZ�ف����)纺+
������*�u39B�x;�n��~�EP��^:�b$qYrp��'kK*�%����z������-�ߵ�p�"��uj�_�~�����t���Mx�w��h����D��gM�U��C2�;�=�Qj!�#V6pL@�l���đ���;�KS;�Ÿ;2Ju�v�ܚ�FϬ��Ν)�E��r��Kw����)3������I�m�S
2����@�z����]wZ��bY�3�qR�7�_���]���(��)l}�%\UD�i�v`��y����#k���kL�0���ُ̹h�"K!Hu�S��{w�T�PA�/�ǩROk*W�ꏡs�'��G�W�Z���f��K������\��A��B��K�^4 ̓u��U�*�M�iɍ�?���4�Ig;��%�H	h!�[�RҠ�%�c���x����X�*�����!#x�l�5�3]���:��J
������I<Id˦�r�
.g�ɸ�T���I`�+��#�J8��	�ņ��{��33�Q��'���M�b]	z�t���J�٘�P���� ?q���( ܍H�o�ښ��H�E��ߚ �	���|�*�a"��[��	��h����>��1Wݿ����,�W�'T����W���c����Uo�C��f�6���< ��w&noȪ�s��i�g�q\Ut����B�h�*��h��ۜ�I숃���!{Y *����3{��J#��a|@�_��B`3@mŧ%w��P��	p�}�z�԰u�S�oK%�;AN�G�z�@�����x���t׽ṋ�dr��l���e�$n�+r4�<N���|�M���<w��k�j
��-w߃���,P{�w��x��Z�0��g�*1��K��u���:>#���\�W�sM�IQ����%�����*���	ZQ����wS�kO�b.p���X����H�e�<�|B�'���q��/��dW�t$"-L�u�7sb�.s���3$M��7��8W���m�-�@(�� �ۭ5XSAH������}ien���
1�t.i{aӚ;��2����T��&����>�=5�'�|��zuK'�^]B+Эߥ�O܉��Pr$w�E�Qk�탷��Nɣ^���izwc�R���NU;}��od^��;�W�������Kd&��`��N �Y2�m,1�l�ɝ�|K
��1�%0wW(��#Cj�l"D5����#XH2�J���������O�ؿ/�>̀�KX��'���\��.f�͈@l�}h��8^"�����b��� �.���h�ǤvZ����{� �)/[�*]��i��J�i�/+��`+�1��=��a��C6��s�ܽJ���;х5^��$�'�Ӯ2
hq�4�OS�ʯ�*T�j�]���k�����Y*�w-�c]-U�"�0m�ۊu�,��r�
9�t���JV|�?!��̆T�˱�Ӡ�e�t����ƕ���ǗL�a�z� �s3�)�o��ˑ���ޜc���~!��:߰8Ϋ���Ŕm����z�!Sv�U�	X�e��j��9�d���ً����2Yo����d^*�}-r��}J�r� +K;N�K�^ё\���()���/4�铔��F�V��܋���	C�tP���:4�������G0��H���X�q;�ӧ{�:��6a�nڵv� �!�l���_�Y�mh�e�II�k��\����lZu"�;:{e�T�Ƽ�d�R��܃~d����M׾ׇ8��I��2K�h�.}4�U�Z8�I����$�D�Y�PfL~�.����CI�S�ILgw��ʚ�e�n#��n�,�z��S��j`��y���GS�ȝ����'�B0�T��C��KW1J�CPY0.e_�a
�{�V��'��*_���J���IE�wN�C�����) ��y2�%p�;�kR#{�S+�r��YQ�Z�Z�?A�,P�}�Q�y!`��ĩ�g���7��A��hq�>a�;"���߮-�����<��ЀQ?I���p�g��p�α�Opj�Qz��e1��U��-������@iy����3�e9Xʿ��5jf�4�J�C"�8�s�(s��-9T��-��[QcI��nYp�x�݀�k�>�|gQ���G��nm��=1yɭ�KOQ5�� �MX)K_|����Up9�{j�$��CQ�(��<��R@z��/���b�)�9h	I����BW���T�F��F侮E&4z�����%У�5�� /.��f�v}F=�Aj?��FlS��P��(G��@E����"¶��)���07��$"~O��i�V;�,y.oj<�"`��un����&.��4�#�o��U����&�S����9�j��$����LX��cٳN\�L�9H�!>�}���hi牳���	���k�Mu
��oFIit�\0�?�k��
�����Pd������5*��Ҩ�,Ё��. W &V��%S����61�uό��"��%��f���"卓7x+~���i��7m�$�y��at��\H��Y5t�E��	7T�@�o:�lbC9��|���[��up6g[�"3@YI�o�6������UL�^���������kj1�d�["�)�`�=��/��NT>�r�D)-m��c��R�Y*�2��>/��}���i#Q�L����Z�%Z�3Ż�~��(������;�����o�4�d��w��%�n���~��x9���P;�p0+��Y����"x���8\��K���T��4g�l���-�T[����b�B�UpW���е�a�$0տO����C%����DNqa�)$���?@_�Mf���R��ѕ�揇@'_b�l��V�����sQ����9�mB�H�Gs;���%,�&��DI��oU�9����h�[O�
���?cc�N�_?o-Ͷ�~\��(��-�n��N���Љ�;�J$��sq�b�$c���y�B�a��U��f��
�#"���U�eE="�V7�U�7�d���#<�͛.�oSy0�]Jo3���~���Q�{�1�2x�p����D�F��I*E�c�O0%#����"'�Kjw�44�N7��-ny�(�w�����?�=�E`��CiT��bD�L�|��z�w
$Q��^`�<���~�?uc-�㿜W5������L�=_W�H�s
z�^Y�03Q�xK�;�e�z�T"�*�9�IG4��F��Jq��}e��ン�9*S��~�D�f�@�%=z�xl���M�S7��kyԳO�d�t�k\��`o�dQ�������H)��k��J{��(*dE�FBge��"?i v�� ���Bu�;�1H�B%�<��.���� 'oP�>��rD��R���.��PPLث�J\:��% ��&b�.�vz�@)w\���([K��J�-�|�&z�rɝ��XuS��ha�j�5���|x�x�θ7�{ìo	I!/? �0טM��(6.�k��M��Ч_�ǚA���]��@��~�b��,�����`��:"��ԗ��Fuޛ�WD�8	y�
Ǧ�HM�Ē���㣐t{kU��*?SZ�e
�CUʳb�
��%}���ũ��Rđ�F�m��8GIF�ù�'��uK�������+ǔЌ����S��㳄�C*�4��
\/z
�K��)b9��}W�����J")acRw��㨗��is�,����9�p)�I�`7��/�~��4�lܢ�)�7���^o��3��8��<9�G��[����(d��l�]e���ʻT|<�M�Z���2N9����r3��T�;a�`����xi�JY�s���c~����MK>y�%�2񔿥��B���e���X���T	v�B����;�i�A��S�̒$x׻AHa��B��@��8��~v�a;�('N�B��1����0.���_cg��zq�/��rw~����5��䵑I��U7>[H�Օ�ĨW`T���Ջq�c*1HƼ�'�q��4��+����Ya����I�/�<9�i�e:n� 3�������[F�y��z�1��G@y�H��������}٥��vf�הB��2N�?Ue�V�֢��f���^/�,��HS�%�f̵�vS�����8�a���&��Myȕ�����,�� R��(�5��a�иFe����6���g��#
�RǇDu�WQHs�?���֮��4���)M3��叼�9�JM[���Dɢ��C!*jYC,��Y���־N�$��b��)y���q��ٙ�cu��]wjxqH=f����b;�=���Q�#r��M�W�˄��~��������P�  EÁsX ��ƕq�?8?�߲K���&LhY�����Y��?=�ϴ��}�]�4�g�߀ۺ@m> ��%()�L��i��a�c�126h�Z�Y��:O�RX��v�ڞC�'�TcE��5sD[���%�s�V�d!� z�1�=�%��T�����#> �Et��m��PHR� �Sz8�V%�ݶ�|j�N)#ʻ��|w� (�mfn�;eI�"���8<���o�Tl���~K�Ŧ�OfIL�uЃ�}b�gf|�1�UNG�4����#�Q�+�v���� ��
�}/������J*D�fvGIԋ$R��	�s�2�]>�|j��I�@�l{H�	�Z^��.�Qo0`;!l��o�7���/������#����bLW�ژ+y�*���#�u:��->ڨo�h�pjtF���q��W���N��n\^��Cc	Im��9L��ҕ���X�`��&z�%ӂ�(K�q��q�+�{��LnO��^�A�j��_(��~3�Rh������Y�bS�9V�H�GN��1|Ñ�C�|kd����K@�D�s�I4nV���p�ҟ�d?]/8\q��J�
=��e5�?k��ܢe7_P�����7�(m�����=���Z���=����ɝ�]\�V�.��g0'����rB�+[9[Qr�tF�\<o�f��(K׿L=l���43Y!��rnpb}D��J��$�L��o�y������k�!�]\�_��"~4�D:\/���R"/�'�:�l�'��|�L��S�2Ğ|0���r�b&2���`���ɱ�{�{ݫIFR�OV���m�hG$��b����� ����;B$�k���C�f'r���i)~�/P�
3Iˠ�L��ɏ����[ܪ�y �v�Ɛ*&壴�4�
o�$�'���6�v��Ԝ����Q{�N5����љ$*s�kgUTF0밶d�8rY�O<`�	Ns;f��do����4���S�l�	mf%�&hN��8�W���g����(V#l}�*�+��;E�b�936��}y��)N�x�Pl��AƊ栔fXO���[�.���#i�)D��W[�����z��{U��z��fq�s�J�2>���٧A���M��Ż1�;g�6�����Tp�CBh�����V����J�\�cl˿�N�M ��z��?���Q�e#����Z1��m���+��x��R�e{v�a�I�uZĵ��ފ�wfB,��p%'��TOX��U��8poU*�NN-
qqTH�5���WH� �����L�i%ꎾ�E+ݞ��	����X�׮HI�V�}�Y(��R�ܕ�h�_�ln��5�n��k�i.�K��d1v�#D��y��U��+�%��v���|�fn���ѐ�R\�Kj2i��ӋY}�FXtX*����|s4�>�KH{f������R�������������b��� Я%��/Z��#
%�Fc�R��RL��+���e	6���꒗v�s����ŗ|bĲ}X�z.���y��L�P�%!:��]1[���\mK�J~�p��a:������j7���$��lBʟ�q���/�� ��ԧ����������� X��u<SKY@'ȹ�qQC�5D#�/��)&���V���=c~E��AKR��;�̧��4��N"{_���w��Z���ʝS|�ߑj;������sl#l{��K��S4T��;+HO
AT�n���"!	;fQ��fL�f��T1F��=&X�;���[��`e_�3��â�u�!���RUC�3t|����>W�8��Ka��bR]��>�G���1痂��	���s�C�|�ux��u��龝~tD��l��󭙋_��P�2<���S��Z ÇL�M�>�څ��ͅ`eµ(U�vY���� �ŏvʑ�bx_5^o���.���x���%�]�(��YZ�Q6����ׇN�][̃Ɖ�+5�o�2
BަB��U��S�:�@�+��a6a&t+`i-�����|�6rOө�����<?�0��x����#ණ�67Z��^�gM���ô{��I��S�.�@��E�\�I�������"����r"i�0m���yA�^��~�K�0�9���쿎�)|��/�����HW��7� K��uÑ�֙_�J�wl��q)ЂJ������E��5�:`����ٞ��G�<ۈ<��|���P󲵝�^�����L|�� ��@t���N5���n��c���;UU�TWɍ@�p��$��Y�*]wբ��<n�`��X� ���co��8�J�g[��h<��:l
��˲X��C�a�ǀƩ_��=
�q1zӸcG��hh
ŎK�/!����FF�z�F�xTfXB((����_v�[1��M�r�x\�lh��2��1�Pn� qE"޺�Kg}�͹T�+?��vwj���y�:�Դ�����B�N���%o��G����)��5��;�"���_�w�T�KW���X-����Ʌ��� ���b;����X�P��x�o޻x&�4�̢����#�u��U�O!5�6�����I�G����=����6��8�p��K�B�i��o�KD�kJjpĞ(��-h����&7�/�5���5�M�����1,]��#�M&�lӂ�H��\q~���2��������
Jg �"r�Yw���h:��r��\��	�IH1l��vG������@^��^���{��1��[��:�� �A����'��*?�3a�<ըjw.B@��v��.ӑ4�U "���/Mᗿ�	A�|��a樨����Q��ƭ E��j*ο��M
��V�s�=x]1oSX(����'�3X�S`��ȱ��<�$�{@�nU�Z�^R}M��2Sxe���Q�4����CU!�h>�K�{CA+UC�:v��/��G������܌b+���4�m� �|,�=�{�N�AhS�G�,��ݧ��D��d��وD)��?��̈�a���.��n�D�F���?1�MCB��J�K�qx�����`�������x���#���I2}��>��~�V"�Ö �7Q�-\������	�&d�􄿝 \�Muv�
L���i�4~� �c9Is0� m��f�t���a4��W��B�Ά>,�}��Ev��������I߭A��u��`����O�V��F~N������E5�L�D U�K��B<V2A�,��`ŀ�jo|A�k`�f�%�L�!W��bMQ�)���s�i�}�����:7sA�F�$�F\�5�<���r��w���J�����CT�Nx��^��%%ҟ'>���(�fB�*�B� �y����Y$ �'�_�rijg��L�.��7[���I�>��ĮM��V�.��	lK��.��ű*l=C�ؤ��4�d�p:�㬼yx��8-�� R�������z�i�,�V���A�I��0���+����܋�Sj�^4w�M)K��m���qZe�Ȉ^�E.�:�]/މ�f2Y�Y:ݧěAl=Eކ����$\�-���
SlJa�{�*6	����Ij"�/H��=?�*�d�K�[U{�4{�&򳈖�u�-#�i;���nL��Uq�a5ي;���*��!�8�~l��r�5�h�ɏ[U��� 	])@ �[��8LǠY4E/*�L+�־��pcQ�\����c�����`jߞ%E��
��Y�&�>K��Q�>St����'g>�'
����2�N�3������ݬz�����M�ϳZ���Ѩ���#83�G��[HI��9ǌ	0�s�z��a����QL:�C�O>K?�+X���瘟[C�k��q�xb%��	?��҆��܄�u�[8�e	 ��~�23�uR5)��Q5���vUP���ܔgC��p���L*���TQ�Z3G̻p3�϶���=Z�m�]��'m����s�4�ಀ���z�~�Z!;c����25^�"��j�==J2܅F'If��>�%wM�XC4���4��	��ο.RԠ���h`��� 9�i<�QR�:;���|�r��Oy3!���pD�L��uB�Wc�n=e{67�&�ʒW~K}�H4��zr|êdg>�G�9�;��1}p���	q�[�y���������,��Be�T_I����!`o;�WD�*2!��pYS��dI��a�Ib�m�;Z}�=�>�;�5s6~s=-D�*�|�"�
O���hp�^~�����G�p�s�H��A���ʮ���]�dTB[.Cl3n��~1EP�gO�h�+��d��}�K������F:a<����Mx�ݿ�Ί8%-7����K�Blg"�	M?�Jt���_�E�dR�񴆙n�w�6(���p&����C*6�>0��E0����P��8"����[W=,Q!k�oܯF)�/n�wV�㞊�������C�����vI�gx�`^���I��}������4�]V_�yE_)O� }�D���N��?!W/��`u�:�N�ʻ=Y�h^��.\})�lЀ"�Rn'ƭ�7`����+
�o�}��|�<o��L����M��,�'ʲ[\z��
�M~�YF��B#��u�S�1��m���h��Y�U'4=)b�)W1����H�OPW�|�7��LM�����ς�(V󳣂^��&�qUMӋoU�b�g�gN������4�������w�����`f�B�hB��ѵ�VmE-��8m�C�[j��}�K�`�0�,TYB�Z�ˊCo1>uU�5�����Y$��V
�����c�l�T�ݳT��wnV�ԗ�4��� J*#^��l� [}����r>��(k/ 6���M��ű�~�����jk�h�Xw6t�od�eƒ�w-�� Z^̮TUS��V�T�� �+�N&>��o'�,FiT����(W1��+�APKh|<��(Թk�f�(jdP�x�#9�bx���C��곯��\3�Ĉ���t��A�m?�3�.��C�A��m��k�9��A��(�d
{�@!�э�%Z V+P7��(c�*�ȒO&�;��݈��u�=q�$~�D'���2QU���E&��Cuh�����
�`g&��d�tEK�+D��Ty���Z�R5�J�%��0Gib$b���2N�?|��O���V��w��(wO ��i&Xi����|Zɓ���{l�u'��He�ݷl��J���9]���~l�+���=��tu2x*-����H�T�h�Jݍ��"�D��D�!�d�`�wP0��	�x�p��v|j�H���{$S�0_E��q����!��g��a.h�I	M׶u:�%�����KXdE{K������/����+��l�W��t˴G~9���ckk���m	�:�۾1U[�"�� ��=�(�>�4G"��F��D�%Z9F*���y{k�Bʐ��5��hX���>9bcй8l�Ξ�Ƿ�w!�eY4�\5\�)�4�C�h��\G���[	ө�M���G&
�ADJ�����D���3�c��|����[�oD�qDQȮaN���μ���_zmK#tM>���2#�摔�%�������)�[�3\C�*�z͈��K��U�Ѫ�	ކ���|�Cy�����o��N
6�k��{�@��:�J��	���p�s�k,����� �%���Y*�wt�0 ����(��3{���й:�3&x������_W�`��,�"|��%XR�*%C��P��[ݯOH��?x }�����D��\P%s�E���ly� n�v
���"�|��z�z8� ��~�K3mи�ƨװ�I�((K��af���-�Wǿ���kkQ�pQ��"�zz��ߧ�)�{p����8��p�Np��^��D�����%�M�CFݽ*��ã�,f��EAB
��$�O�ܔcV=�ՙ�$§��j���	U�[����0��7��h�MK��yĪB�P���;p�4�#nW��!X�\��jX�"� "H�h%y.�S��][ �a���/7�|o95��ng�1~��:�<������]4��m���3g�E��D^��ۉ=C��?��u�� Lb9�7�-�W$-����z�hj�K����ma�A��p�70��� ƨ-���76o`р&�:�(���P�φ8Ɍ��T�Y7����9a��s�gb�}S�l���P��`H]����8�6�\�U:9$@��ѫ��>�򁆀ߺs~kIe�30�E��ǝԝ����f��;*����P�s����04bc��4��kJT;Gm?M~�*��x*��Yժv,���Z&8v�W�j���P�bX�W�0oz�US��1Hb*$��8�n�7�J�~� ��>���V��Ĝ��K���������r���C6��������0�]����]W���m�X6 xfW�!�1$�����%�ƁZ��WH@�n	ߡ ��Jw�~������֚\=�>�M�
�J���������F{�ש�bs!�<X�o�f{z�9b-zL�X�s�V���~��S�����rX�.s?L�ܩ����K�ni�d?��y۾([^uTt	�HݷCq����t0�?Klse�!���-��ɺ���N�bU���=�̆|��C1��P.�ٛש�r�^�9���)�
&DO* o��+ ����d������,�#��:]! ���O|��n}b�q�O!��h0}�����%��|��Fܫ}��edħ���h����q`j�d
�e���+Y��{�Bg4�-t�P�ް�����#��C�?\Е|L��0�jʙd���Ɣ��u�d�����ؓ�W!�ͱ�/���}W^�'�w�;Rt���� ��K�b7)Kũ�E�5��6%-T^��#+��¢d��#5�ҴmSO��(;���%+ aѪh#���M��e�ZZ��מ�[4�w��ae���\�;��A���719�bas�l�����i���:�.i9��b�o��aO�#�p�Rr��-<كкc:#9
��ǃ�0�ɩڹ�$:(��;_v�d#��P JSE��/ �Psb#�����4�%;��%����nJ:X�B�Z�C���/�oیt��Ǯ.pK���b�*�9�gu������U���^�K���h�+vM�!*
W~RH�)q��I�� ��E٬��(��g^��Z��X� /h�]�Z��t�C:ʘq{®)�)��'����RN��f�d}�eq�Q�`/x�-�p͵������p��N����Ie�ڞZ�=��V��U�U�غ6|�V{l�B��?��^��?F���A�lB�ňdu�� }�~�;\ \he2[5�}'N�?��)s�5���&%Ҩ�mq���H��3���vd���s�RL��[�z-�XK1��@eS�ScŢ�[���ra� ���p���T0�7)��r�y�ĥ�V�̙��t�-=C�B���^^ﳸ�,���Vy��!�w��l��<�!Sl�\�Z>�޹����Cu�0ޙ�_�|��0�1�ɫN&����_�HP&��ύ,��߈5�7:��6�vo�'�u.�r4���_���&#�IM������].���׎���p�_}?��"�� �NV?i� �o��U���gA[�Cn�S<j�[�=)b��j�/����g�<�~G�������Ֆ2l�&��r<7�ݽI�{_�!�Y��d��ي�歎_��N^^�r9/�k�D�xuEד���c7vӚ���@�#*�i[ŝ+/�2��L��6;A�C�/�8��G!��"���/��,�5�@�ݚ�2\t��%�x�Kw�gB����z]q�jj�Z^���6�hʀg�fz�N�Q�Lx��M�w�kU��.:�Z� 'c(+S�8
l�w��U�9�cڏ�4[;|�*��&��&��U��d�z�U���޲Ҟ4�Zj$��c��9@��,x�7v�χǞ��גO"`�v́�i��[2��U�MwJ��V1E�v��9&D�Þ������I�d�ا�vz O�P��#�����c��a]�jsBYŰ�ذ��K�����5	7c|w	>n���i����`x�v��T�zP���<��J���[ev�ܹr����m.0���e��o���Yi0^�o|��������+����0"Y��I���׆���BV�G���*
�,�!,�3O�ssfT��[f�x�>J�4x$���}�b��zɅO%�	�ϣq��-��3����tq��~p�e���������`��~#���&d[5bҽ�O�	��6����x���O�KZ�(���7?����L��9�~��#i���BJ��<'G��n��e=��#���\�|�`�Nt�o>)�ɒ�{�q?�NA��#�1*Kj��\Q���-�RTRn��v�B!È�T%�,�^�%'�5o0X_jg2�Y��k�P�U��G�xL@���ޫ��)B�6}�����~��M��,�ݍ!җ����!4��9��g$׶��pmy�G�v��a'~��BbM�\��<+��jw8V��ق-�$��z�W��{���f�V���H腖�����ꯙw��G���ɹTPNRX�N#����l��c�$�A��O��N���Y�#������b�+O
}���J��ۢ~X��֤���,�B4�	}`-���0/i~'hO�\�#�3�U��Zs�� �!�T�C�?�:hizdvC�}�}c�B�'��p3ř���u�[Q�:���'�/�.�I�U4)L\��7�I����F������o�����L�8&q�X�$�� �oG��o����7i���E�F��QY^Pq
'�ύ1�I�"z��	�t���b��o�"���R�(�����=�&���2"��I���z#�c7���g�h��!~~M�K�p�8��~4��*{j�޶���9�o��S�,��W���ș�!|j>�<��{�q���k�I�x.��&��6
�j���X�ٔ�5/������=�7�y����ΰ�U��i��E�}�R�
1��.�om��5t�å��t��:zx?u�m8�<M���������u�-�+� ���`��/"��d�2%�r�='�N�mWz'[���J��NJ��"��ƚ{K�FĈ�#���f0VD������d��u!����	����ԗ0t(VD�G꒸0W~��D���N���d	?)p� �Sک� ���\�c��Vis&S����r�E.ma.��4{7Y\?|v��r�~Xu�/����0����Q^kQ���T/	�������}BZĺȵy���6,��������u�5ȣ���&{��!�;�p�6��m��@K�3L��G���ށ����PA��~{mW��_�'�Q��'_M��4�m�G�{��T@���<i�b�6�ga ?ia�U�
���N�;aJ���tCE���6��s�[=ͣ�GN����`�I(1�x��ej�l焬�˗�i���ߺ��[`{I�x��tE�c��7�4�՟�M���\����)�@S,]�O\���&�!Is`�v�e�(H�U�3WB�Ӄ�S����{�c�o��b�BS�<ҏg�bF]��.�҂4�����Zߗȱ �l���#es�}5պ*܁����6v�0iey���Ĵd u�#f�h՝��vN<�Z)�k���^� ��e��}��Q�j7�n�k%!^\�c���.�"�� ��P�3��x[!X��q�9�(z���{:�J���L��끩G����`��^n෡t;����v��1�FU5��E���7�K��K��P.D�$K#�T����ז������r�a'u�~��򙽜�BHM��p��O���ݔ!�~N�kS�k}��<��9����tjO���ӊB���:n��VTƿ�č��y>��sYfjA
�염|6�3#4^t>��ߙU������G�w��P��!��1�8�cZ*�g��H{�n:α[J݂�2�PN��	!��u/��}�c,�V�'��I��E��k�9��Gx����)z�K�4n�!����	�ܶ�(O
�^B�e^-<F=��T=��*y�j%h#Ki��N���8��GM@H��m����T2s��L�hg�PN���>��'5=���@:�?7:�Z��2���Qv�S�� _�k}��e^%�~!���!~������=����P}��1��ٖ��}aJ((Fw�r�yn�j#�V��'���$��1���o�u���p�g*W���9~�s35=��G�����-	h�f��*�����lj�Q�Yc�@��À�����W�#梬��;mvfl.e��~Λ)c���Gz�F1��#��q\�!��
]��ǟ��y����k�-�?�r��\��Ȏ{���o��4�O	�aa6�1�I�zϤ��)/�!t�s�\CRy�(�e��$/l#�SG���a��T�KOy#+�<3���eD�>��z^Y���R��=���P��ңMJ/A��5��\ ��!IE�y�g*��[��IR�CKX���p�Iи�-[��@C�PO�[���$ ����rW�M~(��&��ɤ�dm��.���,����j4��/&� iM	�ʚƟ}�S��8F��e4�7h9J�&�i�g[Jb.K�X�
�6��nX1�0r� 5Z��J�_2X�6 �hI�x�����.�}�Xg�[���y/o���,j93h��)�a
F�?&P��o��J-u}z89.r����?��jğw��7lf3�	�}�OLf�w9���W0gnX���-����x	p� �T�)�e�ز��~���H-;�u^�`0z��ǌnDA�-	J�I$dAH削@�z����J�]�cI�SO��?�X�G����YP>�B񴒓P��O�~�����M��a@H��3����F���";�k�ڲc��I{t� ���֚)ecPv��J���·4�;&�N跁��4~�S�?�WqpO� ��r1�>�n���T������
S��|��]l�`��MX_�Fh	�3&d�S��D�"��>
��.�� Fi,v�����s�$��1k��a���p�o`*W�Đ��O�c����嶨GL��Z	�t�����vX��4�6�":Q?�ʖ����q����6�S��h��𼚶��e��/
�q�MD���5��l�E�����`XR_�I{��:f�k��Q!=�`�)�d�v��Y��ώ5>���^@f��=�!�?��P�����$����$���.�"�����́�"�W��E�P�MS0�RYd���l�1� de��{�;���D#Z&�Z����q�p���3��ɢ��j� �PUة���c��+��<Fm�5�vy��C���q���Iׂ���#n|��
{�i�ŕ��&ڽ�d,@�n�7ƨKu���*�,��D7��S��zo`���v�	�5��V�ɷ����:	�de_��j��(&WA	m�ƅ*?E�piJ�t�'��B�����9�|�	�&�=��v߁�� j��
�ȀvM)hxr�����\B�gi~�Y[g!� ��/��l�/W�-C)uo�F-�U>ϟ|��5ʽ�@�)�������.�j17�=kZX�l�U�w��&ڸFz�>'F�S��:L�=�'[��}QT� �&���a��~�G���̧��Gٱ|����M+5����W�;�Wr�B�P��Б�Қ�o� i���)~X+����d��o~eo��Yf�-~�trNq��2���>�5��qK��E*�̆
�\�*�y-hZ!a�Ƙ4���DT�hw8S�:���HE#�ꭚ�9?4Jx���a1�����s�����!݈;���c|�7�ϝ��ɿ4�
hq���ND
�`o�f�Ȑ���l�Q�ѱ��M�s5��^޶~�#Z�:;1�`��q��\of}�	�U���c__�P���_���ӽkZ���>A[�PY�b/r��Q���P7���'��}
 K����+�&�\�tY��o��B|OE��v�*~���J 0eZl�%��<�w���` LoW�+��:������d4��i�#p���3q��ZP������m�w����;����3���n���S�qz헦[)j��bܹ1 
���bJZ���� � L)
^5��ܖm{�x����r
U��7��п�s%�n�Kǘ���ӌ�W�+-�9�Ll�Ew)��c�����ܡd3��v�6�������Χ�#6�v���s��m���]�@�x��rFP7ȲL��OD
h:�D<�(e���v��!ejS��L��.
���dZ1{�M�>����2vʈ�\"����?�k�lr!�!�y�h=O�ZV�%��n͋QX:5T�z_{�iK�X���Z�z+ͷծE���`��3B�`D��
�[	k?� "� �W�sЮ�����j�qW
܋hl��"�d���q�Z��6�s�+S��63o	�GƊ:o�p��.��; i��'n�k� j��pU��؞�j�]��U�66�|v&�X���&g/��]�cc�՜�����{=&̶,f/���s��0Z��V18B�t���ȥ(('C� ��<�;+���c΀�a3��'m��_�j�"��v�%f�L�����͘�K�N(?v���I�~?���͗h>�ܪ���f
v�6��������+�7=�o�H��|�f��h]8�wB�G��]�7@`V}�mu���r`��%�F³j��T��7�\����]�mt�V6G3�2�Da�s���e
�|�a��C�M��C�Zt�5k�WD�Z����p����!�:�W�t�B6޹��V�W�V�z�y��F���s�	t�;tb��I�5�8m�;B3��<5�*K&��CWs �mY�J��(���t�4��y�.-4�B��������Ɣ'|����U_2�q-xD�s��f���xT�4m��6���1
:<���T	�:�� >�i��УD�-U��0=���؂�:��vrH��,�<�y�[��YB�lSߣ�CQ�b�����^h?��3��9�{�=�Kb��Ԧ�A�o�����z܂��	���+1�}`�n1�=TicD��e������"��GUM�O�TT�r	��#�<!����j��I�]r/O�Y՜��e����3$GQ]�Q;Э:�U��4��1Q\z[r�xYT�����]���V�k�o�*Q��.Q��,�]�Hz��G2_:F��(���ɷk�e+q�@���BE6���V+�yOu�79���o��;}�'O�\M���/T��pp�q�����P`Y��H1��x����yy��0Ő���2���\�91�p��8�h7$X�R����-�qR}�w劀u2���i�����Zɿ�h�?�y�����e8)J�I��7����"��)I�h��J��{v�K�a�0+�ԯ懋�c�GLq���|H�s�Ӻ�?�I-�ӹ�h�~�/��z���0�6|ngG�w^_֙��GW�ЮP�JZ���v��E����ȳ�xz}��<�N'�Ṷb-ؚ�rg/�������fux��w�?l<��]ÕD�C�QŜ14��Gin�q���1�f�Ve��.֫n�̧/�,�J'/�S�p*�]&��、;}�7tUon���M�p^v�����ˍ�x��3��c.Yp�9����q{��Lv#��
�ߋ1)b_F^1���n���*�Q M���H핁6��R}-5�RX,��7��'�$C�׫p�����~K�JR��h囜h�����\�;�����*�4W���0O\��t��*��e]qAt�K���JX�5��)��z�E�������Y�Dv�/o\��;i�_t����}�px���M�^{e �í�>�?�`>l���g��6Jz�,=MXe_[:���a٧o���.Q���̛����V����4�t9ѩ��P�I�=��N�f���s��$��|�߁�0�~4���0�J���S�ͧY$���5�{%�_��+Z�m$��'�_�sm��1��7��*|!ϳ`b/�v�q)�*�i�?P��/7��u(\��7R�}>��W�`�������un��2&zg�{(�b���80�'��~.�d;,���Ѡ
(�պ����3���&U@T����O��JQ�L�Lx& �U>�}���a}b&����'b]��x���qet�[�OE��1a����qFѕ-U�J-�eJ��E���9v�qH��U#ΔHc�hrc��\oG�t'f<�K�e �s��O��f��r������k�C�����͉?d8_!�|�Ӭc�ɂ^��ڗ��]�ɡ<��}Q�uIɥঞ{3��������^e�X��#�r���|�JcKP�|�D<aߪ�A�����(�C�B�V>��J�g�U�sP��*z���K.L�%��@��0��+i���sEh�nU���~#��Kyl�ox)���>,�I0=��~����,�-�oR���w�_�^7�u�2&�+�مę��6�J��-.��p�p�G!c�j��p�_�6��!4�W%�=]U'c��.��+?�B��Xg��b���a��=��)	���8�Q�޵FZ��D�Jy%pXLY��.�H�P�XQ��#g1���u�l���fS�(�H�e4�Qe6�k�i�����{��G+�A������Q�j��	�����V��i�:�Z��Ғ���})�X��vE8Ѐ��
f;,���\��'��9Hȏ�����h&�˿�ke��H�+��=	 ?��~N�
���s���R������;�jG���8T��ݹu"6?��� y�b�\�;*�g�:�W�y��Cz����"r�Pu���S@�q[���)��F�7������a��)�~�� >�^����H�'(��@�����_C[�M`<��ҊP�bVP���H�xQoC��BM�����C	{�-�v(�#�P���Ǣ�G�"���'i�R���'0<4D�2'��.�p�,v���<P��7�խ�MSf}���W�싫f��^-�\!�l����!� f?Ƀ��K��޺l �=:�������)�����r��L�<����X���u�
B���Ic��Ħkz�:�SX�1�'4Z�2c�A���-�
��(A7��� 3\>�x��`�{�~Z#ym�-�ľ[Д��7ʏ�0��xL}a�V�>��Lt��bi�������yE�=�n��Y=w�%�&D�8a]ǆ�j2X�Y��d`K�ɨ��h�&��~��ˡ)�l�� B{� �mxd�;�qL��|[(��6J�$� �;�Z��:1�ֳd��m[�H��>�Ĩ����:����ۓGd�/�����K��-=���� kmA�H
��-�Ɖ-��^:�~Aoݐ�o.����r��k�L������RA�����s��^�#Q����7�ޞ;�\}U��G�kiJh�ar;|��%�B��D��/䍠��E�J���q�4��M�iy�C�M�L9�~�@3�y��ٺ?����뭨�~��H4&%V�:�!��3�K�S���sDj�Ŭ�12�~�'0�d�غi�"<�ڤ�7\P��2&��Gp�$H�=p���/��=��E.�T�Z"h����Nڝq�� G'�W�8-d�����3*��OO>��"���h�X����M���ev?�+9`4�r�Ծ��7����dsR��zb;aW!������џD9a7�t�m��5|�������A�XU�ص��Zy�z�H�Vj���e�T�:��Jl�l+�0�]7Q�l��?xd|��x�uԡ�iԚ���*'�D*vM���9���j�2J���и�Nñ�UU5A�[�J��M�L���aۻ+a�޾
���$�,�\[��I�W�̴w�w1��,tM;�\�����U��Q	�����m�2}3c�0�b�Sn�R�M.7�����T�<}0�er�k�g���Pǘ-cv��z�������Qq�A^������|>�#���u�[�a#zH	@5= 5a+��l��0����d�9@����b���ȷ��|x����J��&l��t�O��f���`���=��gidâs7�K����Q"����Z?��[a@t̓�!��F���P�V��cs�'��7wچ��%"uv#�p�Eqkq�{^�NIiqD=�ly���>�C��YB33eaa�ɠR�;�8�x�6�Bއ�ZTe�����Cf�(�s��D��:0�+mO�ɭ9B'(��*��� ��XC�Z�[�r�Z������	):J�<,��R����j��>J��Rp�Gc�Ub�f����@H�#�\0Q� ׀�W|������6^n{�/��Ŏ�QnZ�9���-�uV;�o�}k�i:U�|K�c�m�w0Lډ�G���o���b1>�\��-l���䏆�.���B;B���I�=��lyb3Ō�}�Y&k�L�
s���Ǩj��}=�4�s]�kr��i���Vy�̵g�o�0���?��$EcE��Fk�a�J^��kD谱�&8�<ꗶ�bҝЬ�%��Iii�&��W(4sm]C3��J�A�r4N���xsuӈ�\���(�����N�g�GzRvd����˓��7|��`���m��t�������;�v�U|�N�rH1-͙�D��+�$�g�е&�_G���b)=P!iB���� &�"���,����?[�OP��:�+��R�W1� xă!���W����-T^��]�2�OI/� ����J����	���E��OmlMwL�t℣��f�$����[���"%�&4|O����\�����ݖ��/�~.+HX4p�󑫈�u6Ğ�4�w�s�B�ES5�P�i��-����_fۊ*_*��F��%.R����R#�&P>��"�G�!��]�e���<�B��j�~x�z{��Q���x�Ba�[nE>y�U���;ʺ�hV@��4�
<b+^��d�C��t}�WȖ V�&�rk>�� ��ջ�>���R�VAUղ��~�h���7�G��D��5Շ(6b{cP�7脮d��򉃅�%�����������K@����[ǷƉ����yVD�.�5�^AR3m�E��^ ��=��W�����B�3C���қ`蓞	�n���of{EwluT���lңl��0�-��2?q�劽OrxI�B^�By1��zci���K�ŭ̄���U�*}l^W����x�O����������ǡ3>�qg����ڗ=C�2��Tq���&s��.71�9���#Õ�(c�/ X�����߭0��+T�-�tS�jM�n�6�N�46=����\�F��J���a}S���D���V¯i�Έma>���C��Q>��\7)(n�c���Z) �2"�L�@����{&`�D��i��[�#H�l�}U���?SkC$�=���6�A288�)�I�Fn%����:sU�P�T[�&l{�Y����"�p�&Q��O+�ҥ��8y�I��zyȶQ�#������#�&O���(-F&is�8�r-�����q���%�x�{?��06�|TW8�hY1���B�(��+	��^¢N��1z8��XnjefR��\iS

>/,I3�tk}�\�*�^�*�2׶�\B�N�;���b�"U�3��A�%���-��7JF���r�����x�h-��s�%7��n��ew���+߳/�k��w��F��3�0$�H��+ǏS��,?(?�vP�P��5��w����6l��:�J�����jǰ���Z�u�&2�)���jY�IYtH�")���3��I@����nV�
Y>#,��L�!��F�P�^b^����3�����y�I>c��I�h��;�o�߸�Y$=�l�}s�4�XN.̗��3r[�I���;¼37������eN!7����m�9ϒ�/<~���:�e�U��I�w:��n�^�+m�V�e2p����"hH����*r�0T���tݞ��צ�̣ͪ<Ԛ��	)��S��#�P�7:Pz1�
8=p*x�en���OL~J3L8pCN����pHP7�s�NF�f���Z��+���uw�p�s���j6_���M���6��qT�_���E�Z��zQ�Ks�x�������%�WU��M�r�q��h*�t�k�g)��
F����Q��.�n'��6�p�sš}NIR	8���M�SE�ݳ�B��~蜦�b��4R�Y����(}?��:��~�XT�� �����8nJ�m���&Ѓ�/�6��Ҏ���(�N���#�Q$��Vi�����-��f����"���G}��nĎ���V	���a7�����9iJ�������ߍ�-�Ns�@Bja����7�;U�ы\�QҐ��)�O�2U��W���j8[7���ҡ��~��m��d�W��`�;v'}��c8��"�*� .�3�9�鈡�M���]s�v�19I£��`xzk5�_���_oE�k�`JW5#��rϽ2�̛E	�r�|$����ufc㎒x5���+��5+��wQ�A,����ro���mf4�J<���Vԋ�z[ak���s�ߧ�M�;���t����d��,|fM8�$�Lc��ʮ0���֚J�'�yIŝ�t�����Et��bγePM
�cm��pYZb΅̎�u{o룤z��?}^&�����5�������$l�~�ۊ��]h���i�ͬji.~�6{}��o�ڣ2�V��k��Z��
��� ��ûE��)�̮U���|�Gě�ߞ�?�V4P���h5P���� ��x唫�?�AC��K3��̚�G�(�G��t�����ܕ'��K�^)#k:�=�#86�5af
�T:���dY?��B,ӹ߲�X�^cS�%�2��DXZN� X���������lW��i"q٠s>Ԝ>�<�� ���٭�A���^�z�	��t�}2�{�y�vj���^܉�$4-X5|��c,���_P�)'Ɉ�>?u?SB�"\6(6%[���l@=�~�[V�cj
!�Ga2/�Hߤb��0��3� K*��,�����P�cپ��z�x��(4Q��x��V	8Tda�}��ѾKX�F�16x���h��q�n��	�|�4��v�R�4ë�2���,���2�;�ȔOSK�i��I'�r�d1v#���	��V�YEq��d��l��1�R��5��~ArGq3���MS�{2Y�'a�1�"�"�/n�r�Q���g�����K*f,�r�����-�~���0��/#�:��
�G�̈�kz���4��4����b�.GCM�h�o�sn��)���ۖi,Os0Jg(�`�6���0�9�W��c��:|�]�������u��3�T%�~��L.텒|��@��p�Fx��iX��un�D�}�#r�hk��#z����ٔ2�&��O��+h��m�N�T�ZYVZ�w\�ZQ����l?{���/��em�I�0��+rJ�w�9K+뛇P�|b�#�b�| f�;J�4��_0Y��mH9�,�vT��n�����F���y��=��D��^d'Ph�޳�x<9u,U�8�n2������<����WG��Is7���hb,~9�ee�X��k�b'*U�����	��r�Y�n�C��o�9��Uڝ��9q@G��6k��q�;��G*�Y������b����F(IUj/(t6xJ��ؤ}���B�k~��f��6�&�T��������aW�S��V	N�b�/�Ǥ�,L��!] �����������9D!]$1Z��j�B��_��:�L�b��Yxa?Q���P��߂,���is;)!<���`�y�#Z�p���+,��a@�\�u�x�N���6]��K��*_��^S69�މ�#?�@��G�5DLj|w`l*�[%?	�\z8�E�{R�e�)o`��	�ns��jB�ƕ��T@�RpF;�����P��O����H`��Y��h�9��6 �.���J��{�܍#Y>�Q�����%xCF���p!C'�Y6W���@��zR���*e�����ʢ����4]K��E������L�
O�3����\�ҷ�;U5���n)�xx ���GIHp)�/}�D�`J�bne�Xe~ۑ�3���u�����͸��)՚�uڍEd�tY-����+`�����߉������6/m�ˌ�ε[)l-�<��"�Կe�x�F`֠sS�x네i�Ko �60�6�j����#���@u"�g�e�0c�uT���R�.�O6���gv�=�R� &Xۘ�>���'"�� �K:��.�h&�F���W�0j��Q�����I\�ٌ{�p��XV}&�����:�8��Cp	����Rш�K���\�J�M�N0 ck8��|5�RV��c�9H�p���=ù(�צ����b�����^Q���c8�Ym�u���d+�y`=+���@�Z8��R硫I^1���1�m�曋-B1Q�x��a�6D��0�������tn d��͙Y���8g�)*��H�o��b(tO[ P�
Ш���Y>����Z�b!�KؒR� r���k��_{�ĺ����Ye�ƍI9z5�_EPv_��P�J�I�I�C`�}��6L Ÿr���e�Qg�&���
����PD�5og>7����I���J(˹/Q�IR�"ϼ��>��?ñI6�M�zB�@��'�n�ԅj��}�Τ��\�>����u�������,��R�?�f��z�dfʻ��b�3��p0��S�Qw�R m��2��4ZpR'�ÐcQi#ǃZe�]��<Bتf~��%(+�i��|=�5x�鷨�?�'V��!�}v�Y_�I]ծ����_rL'm��Lj�U�cyGV-^妘�$���B�µ�.��0a��U���Q���'�or԰6�h�Z�~~�
��8�@}�x�}u��t��T�&�s�:wAn��q�)�-i�^-#P�D�
�+P�j����>&}�V��4�n��/�d.W]�������ee.�����O6�����"f��cgԴ�Y��<.�ĺ܇�̔|���4���Xc6�Lyp��������睰,�	1^�R��f�A�������L���Z�|U���}a�
~�冂!9��6Pꞟh������������f{b����v�c#��m�uo����S���#���]Ɵ-��Ʉ�0-�x���T���F��TWn�����r�nvS�}�#I�;��u� �����b��6(��܊@'���%KO���8�R^��+͗,�4\���i0�i�:�s�`�N��R²RY5�>x�L�����{�q�����HX�J$(|�*{�[��\����(>�o2�M���
�P����ɳYm�v�����=��h��t�,`Q�����
$��`����W˚��Ǜ��2̍9�/o��㊲�ue]٣�m�gks��jG�tVƗ��͐�,��7UnQ��2R��	�@�Z��uY&�v�"2 �t
"�ղ�P�3\e�f��W"S��#@��i0!�������F�MÕ�������D�tX:׌S�
mְ#��ŵy� �{<^���C/��h���ыp9��$�S6��R_�,�,w�W��<�e�.ly��|r�����L�녩_������#��\�֬�fCxz�\GRj��u[s�<��:��� FS�ݎ<���K�+��E~�*q�BXsno-/P255�|̆�S�8Oe&uC�#��"Y����ѽ�G}�gxY��8���J=��㷰���.�7�qqN�f���w<YӜq��6DK�#�q����Ub	$���ŵ�_U�\��1�'�[�WO�5ѝ\���,�s��N�ֆӚ�l�k��l&��2�Xtb�<r���\[j%�Q��پ�7�H$+>i�΢�ʞ��s���'�����B��"���@��J��e�d<�`)�Ù�F� rب �;W�c:F%��_���^��9e�CN"��l˵�p�5���O���H�Z��:�Y��`U*��F7�$�	�}��P����_��8�`JE���ս�p�k��-���iN�M�����;G�se��_Ãty�"�o��H����ʰ8��p�a'�qO�N�Y��˙�փTC���p3'(�9	�\x�Si�C��gǲ��&���τW̅t����5��Ĵy�ta?������9�z�W^�9���W�����j�Vܹ5����6E�ł��6k>���B[q�,��񐧆q��l�"+����h��b����jb�h
��	��s�����OS!�Φ[hƻׇy9��쫒����c|�X�}3y��\/��p�l�ZVc��Z��+�K��N�b�,�*^$9����>��h���'�֥�b��*� ��.s	'83��	���x���*����ڑWS	�Z��ۍ ��(u�g%'9�
K�%�'��4ugz��`��3���%$>��As�ڛ��\ٳ�c"�?F��K�v��K���"��X�����}��¾T�����l1��a�%���U8f�u^��W������b���)��2�TK��9���;�U���x)�S��������"���N��)�dVv��V�'J5+��h��U#�+LWr�٘"�����R�ҟ\�D�6���w���� ӻP����yu(NE����oY1_��`j-�dN��tal��r �?n�E�Y|�{�[]J.c��4z ��~e#���"V�ZU)����c�J���_D���D�,���A��,���Z:稛I����s����^�!y�[�D�GΠ��7E�Us��q�Z��@�S���8��/K@E��ʲ�,=�3P^ ����p�xy�������i�0!�
Cԉ��x��u
Q�L�2 ��qSGg��kb.˴�Cy0�KV𭂁Z�*����W�2�^�	��i�!�gE@�jI;b����+n@׃�F��'Qx�Ȟb��R�m	�䋎�AW����f�欼��,�0�	����ZT"��ADŞ+(���]+�g�bXلs���8�� �1O:+�T����(��i�>��#��s�\�nU=}����;���t��֧�G�н��p�q�| �Adp��{q�i 6+��2Ԉ�?h|����+T�n�W�4`,,t���Zĝ���R3���sm�� ����*ߤ��c��xX�3ՄJ��� �A����0VQ��v�=9vRE�i�(�B� ,�SMc~�H���zX6N���S��������Ә�c`���QG<�����VQ�d�,�q�n5�y:�=y��[%񽄱36�0D�1�D��ܜ�S��5�K:6r*���Jk��"��>\Ķb�\y�����E4��#X:�0j��z�'����N/1Pd9�J����Fs#�RPN�󛍇L��qkP;���z�g�)��؊-0��D�uQBP� u����Г�0�i�����8�ءVB�����dۅn�E��,�"`�v$��y�mK81�xa$��b'`�P�b�m�b��%���jS
Z�,�@�` ��!�Z/N�&��m�W��|���+8kl���Zu�*�=`��y�cH�����dU~����P[�n3Y�� ��
����.9��	Ca��=
����:Q����	����l�0�׭����4�9����"��.#=�JLOOh&0�UA����)Љ�_����TJ-�L��?�g4���y>ɵ#ۗfz�X:�iA-��x�-Y�&�����Ϙ�����,hv�7A���r�)�
��Mk�l(L��'�Y��e6�6�i�k6�r�*��U/��Cwz���cPWл"y�]��%�i�p��t
'C��J�kkZ�\F����)��;Le<�q��c���A������&!�N���=�[���u3��b���:��m�'
��l7���>m�� ��O���#&��b���f_��8��ky�y�Q��d����G�  �OK�t�)%Q�5�Tb}��&Юi���wv�D$Zm:G�?p�>�Z0J+A���,����Y�'#���"HO�7�(���{L႖t�M�w扴O]X�[��
2��d�6N��a@5�2-��5uu��ۋ]O��9���ET��Zn����3��[����9�sH���aO�4c���>Qz	x���D��qX�k�ܣ_���*]TdY̡�]�B�kT��M�DǙ�� �.�hJc���)�D�'ZNjnt+hE��Q`ς	��ru�fKIy��-��ic�K�5�ApP�����k�RE��-G2Ѓ��ˉz]g]�c�8 m�J�	E5I��3�{�J��]�"k����<���P��1V����?,�A�8��Ď�����OD F1x0�DIJr۲����
Wמ�9��3o�a��u�#���U��W��|?�]-��#H��N�Ó)婬ܣ[��şR���,�p}�@n��ASO�5"bb��}���,��E�p����]	���g�"G�V��ص8�i��ݣ�.�Tg�}� �A�B�1)rc�g#|Ŏ(YQb_z�=����G%־)ղs�_�v˪/��7qH�5W��n�F�@e��H�`r6�{��GSy?���-L��:��qL�����F�n������iM���I�icq���hdR��LZQ\^���:�5���r����L"c����)琜�����.��Ү�9v�)E��҉_.4dOO�j��̗�i7D�Nρ�+����H�C-�>c~"Q���\Mc��ԯ�}��f���*�l�'���&"!��ݣ ʎz����p���7��ণo��z�א�:;�l#��ۃ�a�������z]ļ8� ���ASOu"�Ϭ���2�����5)�h�|Sci���'߅[	���E�p���璻�1O*�ɯ������Ur%��N��fs�B���;�X�y��!���:��駺v?�mױ��9��<��tG�Ê��Jz3��$j��%ԌP�]�:��������be�%m"9�'�{To�3g$1&.ipc�C;O�]alf�ܶ �
I�6
��T�2�KN�XɎ�ȏ�'Qϑ�k���C���t�X���"�4��}�9��U�c�9��[O��q��yY���6Ovf�+|�i'.��<a��8pP\���)|�!؉mвk2��#O�+(�a���eZz�J������`�M4q�����`�1W�4B]�Q�M)��/Gy#�e�r�8uY�u��cN�W�O�l[���tZ(�d����$\۟���g���*�7QA�C���P�eo��R�ǚ�-Lf�-�)�] �l�？�(ǅ�6��i�43W��UA�!�x�P:d+��:=:PC��/�ٻÊ<hX?����{!�l]�i��骂�itb{e�s����E	���9pc��_�٣-��������dUN�~"��:������9d�@�Ɏ�l����P�7�*�U��cY̛�Z�Y=�?���RM�v�0����*���I�:ڝ4�@�5�I�;�
A�Y4o�ed6G�6�"��lu�@��%��.���/�����⢡ѱj��zJԓ���e̷Ҙ��V�7Su	���!J��^�Ҙ�{h붬W�����[�E���w��ˈ�tJ��v�D��Ct��ԍAU�y��M�ݽ}�XH���j�t�ʚ�@E�q�=
���*+'�f��3n$0��@͐K�:u|62g�	}�)��3pKxx$ '��%��z�
1^�ב6�&��8���|`�ϩ������W�n��0w��P�먖Ѡ�ck�BɽHh�VF"�`lM{ܒ�|�V/s'���n900���m�(1B��"4��2i���p�]��6�7|k���~
bЧu{nx��ȯ�>��D��\�.ى�z�	�O٣�z��e���!�a��ȓ����z�`·������t�8)�C*�1L�^����TDg�֝}���0�ĝ=�W/�b�	���&����K����-q���_���[��z=�����.a�E��n��K����g�����1���	���ާPbQ�|e���⍂�	PJK��f�z�5n��Jv�.����3���L�y^t�O�ؔ�x��f����g{���H�&�{�@DQԢ��#�sHEl$]���H���I�XQMʕ�P[�i����>�!(�&�w8V$����  d�?.����YJ�Ռ����	��Y�C������ŪP��b�&�?6��,Jz]+�O��nJ���] H�C� ��$�=�1�����Q��
�mq>>� ��q楕6ؚ����g�2��'��s�Oi��+�)<��ø��l��h��7�2 �@fw�+��v?��K�tK=Y��*�	Z��?�w^������Y8%�2��i"�1�!��a�/]�{r5g�FJѓD�J��Ý�x]C���46 �Z'����G{zI
B���p"�휅��Pl��>n�߉o([ܿ��j!�b��%?Z��Q��
ʸ���I���!�G<}u�J4y��&@����d.��+xNv�;NW7�ȗL쯚�
��Ķe�S%GiN˷�@F�������o����92��H;�